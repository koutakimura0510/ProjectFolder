
//
// Verific Verilog Description of module MTopTi180MIPI25GRxHDMIV101
//

module MTopTi180MIPI25GRxHDMIV101 (MipiDphyRx1_RESET_N, MipiDphyRx1_RST0_N, 
            MipiDphyRx1_STOPSTATE_CLK, MipiDphyRx1_STOPSTATE_LAN0, MipiDphyRx1_STOPSTATE_LAN1, 
            MipiDphyRx1_ERR_ESC_LAN0, MipiDphyRx1_ERR_ESC_LAN1, MipiDphyRx1_ERR_CONTROL_LAN0, 
            MipiDphyRx1_ERR_CONTROL_LAN1, MipiDphyRx1_TX_REQUEST_ESC, MipiDphyRx1_TURN_REQUEST, 
            MipiDphyRx1_FORCE_RX_MODE, MipiDphyRx1_TX_TRIGGER_ESC, MipiDphyRx1_RX_TRIGGER_ESC, 
            MipiDphyRx1_DIRECTION, MipiDphyRx1_ERR_CONTENTION_LP0, MipiDphyRx1_ERR_CONTENTION_LP1, 
            MipiDphyRx1_RX_CLK_ACTIVE_HS, MipiDphyRx1_RX_ACTIVE_HS_LAN0, 
            MipiDphyRx1_RX_ACTIVE_HS_LAN1, MipiDphyRx1_RX_VALID_HS_LAN0, 
            MipiDphyRx1_RX_VALID_HS_LAN1, MipiDphyRx1_RX_SYNC_HS_LAN0, MipiDphyRx1_RX_SYNC_HS_LAN1, 
            MipiDphyRx1_RX_SKEW_CAL_HS_LAN0, MipiDphyRx1_RX_SKEW_CAL_HS_LAN1, 
            MipiDphyRx1_RX_DATA_HS_LAN0, MipiDphyRx1_RX_DATA_HS_LAN1, MipiDphyRx1_ERR_SOT_HS_LAN0, 
            MipiDphyRx1_ERR_SOT_HS_LAN1, MipiDphyRx1_ERR_SOT_SYNC_HS_LAN0, 
            MipiDphyRx1_ERR_SOT_SYNC_HS_LAN1, MipiDphyRx1_RX_LPDT_ESC, MipiDphyRx1_RX_DATA_ESC, 
            MipiDphyRx1_RX_VALID_ESC, MipiDphyRx1_RX_ERR_SYNC_ESC, MipiDphyRx1_TX_LPDT_ESC, 
            MipiDphyRx1_TX_DATA_ESC, MipiDphyRx1_TX_VALID_ESC, MipiDphyRx1_TX_READY_ESC, 
            MipiDphyRx1_TX_ULPS_ESC, MipiDphyRx1_TX_ULPS_EXIT, MipiDphyRx1_RX_ULPS_CLK_NOT, 
            MipiDphyRx1_RX_ULPS_ACTIVE_CLK_NOT, MipiDphyRx1_RX_ULPS_ESC_LAN0, 
            MipiDphyRx1_RX_ULPS_ESC_LAN1, MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN0, 
            MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN1, MipiDphyRx1_WORD_CLKOUT_HS, 
            MipiDphyRx1_LP_CLK, MipiDphyRx1_RX_CLK_ESC_LAN0, MipiDphyRx1_RX_CLK_ESC_LAN1, 
            MipiDphyRx1_TX_CLK_ESC, oAdv7511Vs, oAdv7511Hs, oAdv7511De, 
            oAdv7511Data, iAdv7511Sda, oAdv7511SdaOe, iAdv7511Scl, oAdv7511SclOe, 
            oLed, iPushSw, iSCLK, iBCLK, pll_inst1_LOCKED, pll_inst1_RSTN, 
            iVCLK, pll_inst2_LOCKED, pll_inst2_RSTN, oTestPort, jtag_inst1_TDI, 
            jtag_inst1_TCK, jtag_inst1_TMS, jtag_inst1_TDO, jtag_inst1_SEL, 
            jtag_inst1_DRCK, jtag_inst1_RUNTEST, jtag_inst1_CAPTURE, jtag_inst1_SHIFT, 
            jtag_inst1_UPDATE, jtag_inst1_RESET, jtag_inst2_CAPTURE, jtag_inst2_DRCK, 
            jtag_inst2_RESET, jtag_inst2_RUNTEST, jtag_inst2_SEL, jtag_inst2_SHIFT, 
            jtag_inst2_TCK, jtag_inst2_TDI, jtag_inst2_TMS, jtag_inst2_UPDATE, 
            jtag_inst2_TDO);
    output MipiDphyRx1_RESET_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_RST0_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTROL_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTROL_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_REQUEST_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TURN_REQUEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_FORCE_RX_MODE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [3:0]MipiDphyRx1_TX_TRIGGER_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [3:0]MipiDphyRx1_RX_TRIGGER_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_DIRECTION /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTENTION_LP0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTENTION_LP1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ACTIVE_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ACTIVE_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ACTIVE_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SYNC_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SKEW_CAL_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SKEW_CAL_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_SYNC_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_LPDT_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ERR_SYNC_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_LPDT_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]MipiDphyRx1_TX_DATA_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_VALID_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input MipiDphyRx1_TX_READY_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_ULPS_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_ULPS_EXIT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_CLK_NOT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_CLK_NOT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_WORD_CLKOUT_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_LP_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_CLK_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511Vs /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511Hs /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511De /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [15:0]oAdv7511Data /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iAdv7511Sda /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output oAdv7511SdaOe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iAdv7511Scl /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output oAdv7511SclOe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [5:0]oLed /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [1:0]iPushSw /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iSCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iBCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_inst1_LOCKED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output pll_inst1_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iVCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_inst2_LOCKED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output pll_inst2_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [25:0]oTestPort /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst2_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    
    wire rBRST, rVRST, rnVRST, \la0_probe18[0] , \MCsiRxController/MCsi2Decoder/rHsSt[0] , 
        \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs , \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd , 
        n106, n107, la0_probe15, la0_probe2, la0_probe0, la0_probe16, 
        la0_probe4, la0_probe1, la0_probe8, la0_probe12, la0_probe11, 
        la0_probe7, la0_probe14, \la0_probe5[0] , la0_probe13, \la0_probe6[0] , 
        la0_probe3, la0_probe9, la0_probe17, \MCsiRxController/wHsPixel[0] , 
        \MCsiRxController/MCsi2Decoder/wFtiRvd[0] , wCddFifoFull, n129, 
        n130, \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] , 
        \MCsiRxController/wHsValid , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] , 
        \MCsiRxController/MCsi2Decoder/rHsSt[2] , \MCsiRxController/MCsi2Decoder/rHsSt[1] , 
        \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6] , 
        \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4] , 
        \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2] , 
        \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] , 
        \MCsiRxController/MCsi2Decoder/wFtiEmp[0] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[16] , n183, n184, \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] , 
        \MCsiRxController/wHsPixel[1] , \MCsiRxController/wHsPixel[2] , 
        \MCsiRxController/wHsPixel[3] , \MCsiRxController/wHsPixel[4] , 
        \MCsiRxController/wHsPixel[5] , \MCsiRxController/wHsPixel[6] , 
        \MCsiRxController/wHsPixel[7] , \MCsiRxController/wHsPixel[8] , 
        \MCsiRxController/wHsPixel[9] , \MCsiRxController/wHsPixel[10] , 
        \MCsiRxController/wHsPixel[11] , \MCsiRxController/wHsPixel[12] , 
        \MCsiRxController/wHsPixel[13] , \MCsiRxController/wHsPixel[14] , 
        \MCsiRxController/wHsPixel[15] , \wHsWordCnt[1] , \wHsWordCnt[2] , 
        \wHsWordCnt[3] , \wHsWordCnt[4] , \wHsWordCnt[5] , \wHsWordCnt[6] , 
        \wHsWordCnt[7] , \wHsWordCnt[8] , \wHsWordCnt[9] , \wHsWordCnt[10] , 
        \wHsWordCnt[11] , \wHsWordCnt[12] , \wHsWordCnt[13] , \wHsWordCnt[14] , 
        \wHsWordCnt[15] , \wHsDatatype[2] , \wHsDatatype[3] , \wHsDatatype[4] , 
        \wHsDatatype[5] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1] , 
        \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3] , 
        \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5] , 
        \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] , 
        wVideoVd, n268, n269, \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] , 
        \MCsiRxController/wFtiEmp[0] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] , \wVideoPixel[0] , 
        \wVideoPixel[1] , \wVideoPixel[2] , \wVideoPixel[3] , \wVideoPixel[4] , 
        \wVideoPixel[5] , \wVideoPixel[6] , \wVideoPixel[7] , \wVideoPixel[8] , 
        \wVideoPixel[9] , \wVideoPixel[10] , \wVideoPixel[11] , \wVideoPixel[12] , 
        \wVideoPixel[13] , \wVideoPixel[14] , \wVideoPixel[15] , n304, 
        n305, \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] , 
        \MVideoPostProcess/rVtgRstCnt[0] , \MVideoPostProcess/rVtgRST[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_m_en_1P , \MVideoPostProcess/inst_adv7511_config/r_last_1P , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] , \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P , \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P , 
        \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 , \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] , 
        \MVideoPostProcess/inst_adv7511_config/w_ack , \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] , 
        n386, n387, \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] , 
        \MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] , \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] , 
        n441, n442, \MVideoPostProcess/mVideoTimingGen/rVpos[0] , n444, 
        n445, \MVideoPostProcess/mVideoTimingGen/rFvde[0] , \MVideoPostProcess/mVideoTimingGen/rHpos[0] , 
        \MVideoPostProcess/mVideoTimingGen/dff_41/i4_pre , \MVideoPostProcess/mVideoTimingGen/rVpos[1] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[2] , \MVideoPostProcess/mVideoTimingGen/rVpos[3] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[4] , \MVideoPostProcess/mVideoTimingGen/rVpos[5] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[6] , \MVideoPostProcess/mVideoTimingGen/rVpos[7] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[8] , \MVideoPostProcess/mVideoTimingGen/rVpos[9] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[10] , \MVideoPostProcess/mVideoTimingGen/rVpos[11] , 
        \MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre , \MVideoPostProcess/mVideoTimingGen/rFvde[1] , 
        \MVideoPostProcess/wVgaGenFDe , \MVideoPostProcess/mVideoTimingGen/rHpos[1] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[2] , \MVideoPostProcess/mVideoTimingGen/rHpos[3] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[4] , \MVideoPostProcess/mVideoTimingGen/rHpos[5] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[6] , \MVideoPostProcess/mVideoTimingGen/rHpos[7] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[8] , \MVideoPostProcess/mVideoTimingGen/rHpos[9] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[10] , \MVideoPostProcess/mVideoTimingGen/rHpos[11] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] , wVideofull, 
        n481, n482, \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12] , 
        n508, n509, \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] , 
        n525, n526, \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12] , 
        n552, n553, \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] , 
        n569, n570, \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12] , 
        n596, n597, \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] , 
        n613, n614, \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12] , 
        n640, n641, \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0] , 
        n657, n658, \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12] , 
        n684, n685, \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0] , 
        n701, n702, \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12] , 
        n728, n729, \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0] , 
        n745, n746, \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12] , 
        n772, n773, \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0] , 
        n789, n790, \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12] , 
        n816, n817, \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0] , 
        n833, n834, \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12] , 
        n860, n861, \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0] , 
        n877, n878, \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12] , 
        n904, n905, \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0] , 
        n921, n922, \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12] , 
        n948, n949, \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0] , 
        n965, n966, \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12] , 
        n992, n993, \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0] , 
        n1009, n1010, \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12] , 
        n1036, n1037, \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0] , 
        n1053, n1054, \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12] , 
        n1080, n1081, \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0] , 
        n1097, n1098, \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12] , 
        n1124, n1125, \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0] , 
        n1141, \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12] , 
        n1167, n1168, \MVideoPostProcess/rVtgRstCnt[1] , \MVideoPostProcess/rVtgRstCnt[2] , 
        \MVideoPostProcess/rVtgRstCnt[3] , \MVideoPostProcess/rVtgRstCnt[4] , 
        \MVideoPostProcess/rVtgRstCnt[5] , \MVideoPostProcess/rVtgRstCnt[6] , 
        \MVideoPostProcess/rVtgRstCnt[7] , \MVideoPostProcess/rVtgRstCnt[8] , 
        \MVideoPostProcess/rVtgRstCnt[9] , \MVideoPostProcess/rVtgRstCnt[10] , 
        \MVideoPostProcess/rVtgRST[1] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] , 
        \genblk1.genblk1[0].mPulseGenerator/rSft[0] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] , 
        \genblk1.genblk1[0].mPulseGenerator/rSft[1] , \genblk1.genblk1[0].mPulseGenerator/rSft[2] , 
        \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] , \genblk1.genblk1[1].mPulseGenerator/rSft[0] , 
        \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] , \genblk1.genblk1[1].mPulseGenerator/rSft[1] , 
        \genblk1.genblk1[1].mPulseGenerator/rSft[2] , \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] , 
        \genblk1.genblk1[3].mPulseGenerator/rSft[0] , \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 , 
        \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] , \genblk1.genblk1[3].mPulseGenerator/rSft[1] , 
        \genblk1.genblk1[3].mPulseGenerator/rSft[2] , \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] , 
        \genblk1.genblk1[4].mPulseGenerator/rSft[0] , \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] , 
        \genblk1.genblk1[4].mPulseGenerator/rSft[1] , \genblk1.genblk1[4].mPulseGenerator/rSft[2] , 
        \edb_top_inst/n3116 , \edb_top_inst/la0/la_run_trig , \edb_top_inst/la0/la_trig_pattern[0] , 
        \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig , 
        \edb_top_inst/la0/la_capture_pattern[0] , \edb_top_inst/la0/la_trig_mask[0] , 
        \edb_top_inst/la0/la_num_trigger[0] , \edb_top_inst/la0/la_window_depth[0] , 
        \edb_top_inst/la0/la_soft_reset_in , \edb_top_inst/la0/address_counter[0] , 
        \edb_top_inst/la0/opcode[0] , \edb_top_inst/la0/bit_count[0] , \edb_top_inst/la0/word_count[0] , 
        \edb_top_inst/la0/data_out_shift_reg[0] , \edb_top_inst/la0/module_state[0] , 
        \edb_top_inst/la0/la_resetn_p1 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/la_resetn , \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/internal_register_select[0] , \edb_top_inst/la0/la_trig_pos[0] , 
        \edb_top_inst/la0/la_trig_pattern[1] , \edb_top_inst/la0/la_capture_pattern[1] , 
        \edb_top_inst/la0/la_trig_mask[1] , \edb_top_inst/la0/la_trig_mask[2] , 
        \edb_top_inst/la0/la_trig_mask[3] , \edb_top_inst/la0/la_trig_mask[4] , 
        \edb_top_inst/la0/la_trig_mask[5] , \edb_top_inst/la0/la_trig_mask[6] , 
        \edb_top_inst/la0/la_trig_mask[7] , \edb_top_inst/la0/la_trig_mask[8] , 
        \edb_top_inst/la0/la_trig_mask[9] , \edb_top_inst/la0/la_trig_mask[10] , 
        \edb_top_inst/la0/la_trig_mask[11] , \edb_top_inst/la0/la_trig_mask[12] , 
        \edb_top_inst/la0/la_trig_mask[13] , \edb_top_inst/la0/la_trig_mask[14] , 
        \edb_top_inst/la0/la_trig_mask[15] , \edb_top_inst/la0/la_trig_mask[16] , 
        \edb_top_inst/la0/la_trig_mask[17] , \edb_top_inst/la0/la_trig_mask[18] , 
        \edb_top_inst/la0/la_trig_mask[19] , \edb_top_inst/la0/la_trig_mask[20] , 
        \edb_top_inst/la0/la_trig_mask[21] , \edb_top_inst/la0/la_trig_mask[22] , 
        \edb_top_inst/la0/la_trig_mask[23] , \edb_top_inst/la0/la_trig_mask[24] , 
        \edb_top_inst/la0/la_trig_mask[25] , \edb_top_inst/la0/la_trig_mask[26] , 
        \edb_top_inst/la0/la_trig_mask[27] , \edb_top_inst/la0/la_trig_mask[28] , 
        \edb_top_inst/la0/la_trig_mask[29] , \edb_top_inst/la0/la_trig_mask[30] , 
        \edb_top_inst/la0/la_trig_mask[31] , \edb_top_inst/la0/la_trig_mask[32] , 
        \edb_top_inst/la0/la_trig_mask[33] , \edb_top_inst/la0/la_trig_mask[34] , 
        \edb_top_inst/la0/la_trig_mask[35] , \edb_top_inst/la0/la_trig_mask[36] , 
        \edb_top_inst/la0/la_trig_mask[37] , \edb_top_inst/la0/la_trig_mask[38] , 
        \edb_top_inst/la0/la_trig_mask[39] , \edb_top_inst/la0/la_trig_mask[40] , 
        \edb_top_inst/la0/la_trig_mask[41] , \edb_top_inst/la0/la_trig_mask[42] , 
        \edb_top_inst/la0/la_trig_mask[43] , \edb_top_inst/la0/la_trig_mask[44] , 
        \edb_top_inst/la0/la_trig_mask[45] , \edb_top_inst/la0/la_trig_mask[46] , 
        \edb_top_inst/la0/la_trig_mask[47] , \edb_top_inst/la0/la_trig_mask[48] , 
        \edb_top_inst/la0/la_trig_mask[49] , \edb_top_inst/la0/la_trig_mask[50] , 
        \edb_top_inst/la0/la_trig_mask[51] , \edb_top_inst/la0/la_trig_mask[52] , 
        \edb_top_inst/la0/la_trig_mask[53] , \edb_top_inst/la0/la_trig_mask[54] , 
        \edb_top_inst/la0/la_trig_mask[55] , \edb_top_inst/la0/la_trig_mask[56] , 
        \edb_top_inst/la0/la_trig_mask[57] , \edb_top_inst/la0/la_trig_mask[58] , 
        \edb_top_inst/la0/la_trig_mask[59] , \edb_top_inst/la0/la_trig_mask[60] , 
        \edb_top_inst/la0/la_trig_mask[61] , \edb_top_inst/la0/la_trig_mask[62] , 
        \edb_top_inst/la0/la_trig_mask[63] , \edb_top_inst/la0/la_num_trigger[1] , 
        \edb_top_inst/la0/la_num_trigger[2] , \edb_top_inst/la0/la_num_trigger[3] , 
        \edb_top_inst/la0/la_num_trigger[4] , \edb_top_inst/la0/la_num_trigger[5] , 
        \edb_top_inst/la0/la_num_trigger[6] , \edb_top_inst/la0/la_num_trigger[7] , 
        \edb_top_inst/la0/la_num_trigger[8] , \edb_top_inst/la0/la_num_trigger[9] , 
        \edb_top_inst/la0/la_num_trigger[10] , \edb_top_inst/la0/la_num_trigger[11] , 
        \edb_top_inst/la0/la_num_trigger[12] , \edb_top_inst/la0/la_num_trigger[13] , 
        \edb_top_inst/la0/la_num_trigger[14] , \edb_top_inst/la0/la_num_trigger[15] , 
        \edb_top_inst/la0/la_num_trigger[16] , \edb_top_inst/la0/la_window_depth[1] , 
        \edb_top_inst/la0/la_window_depth[2] , \edb_top_inst/la0/la_window_depth[3] , 
        \edb_top_inst/la0/la_window_depth[4] , \edb_top_inst/la0/address_counter[1] , 
        \edb_top_inst/la0/address_counter[2] , \edb_top_inst/la0/address_counter[3] , 
        \edb_top_inst/la0/address_counter[4] , \edb_top_inst/la0/address_counter[5] , 
        \edb_top_inst/la0/address_counter[6] , \edb_top_inst/la0/address_counter[7] , 
        \edb_top_inst/la0/address_counter[8] , \edb_top_inst/la0/address_counter[9] , 
        \edb_top_inst/la0/address_counter[10] , \edb_top_inst/la0/address_counter[11] , 
        \edb_top_inst/la0/address_counter[12] , \edb_top_inst/la0/address_counter[13] , 
        \edb_top_inst/la0/address_counter[14] , \edb_top_inst/la0/address_counter[15] , 
        \edb_top_inst/la0/address_counter[16] , \edb_top_inst/la0/address_counter[17] , 
        \edb_top_inst/la0/address_counter[18] , \edb_top_inst/la0/address_counter[19] , 
        \edb_top_inst/la0/address_counter[20] , \edb_top_inst/la0/address_counter[21] , 
        \edb_top_inst/la0/address_counter[22] , \edb_top_inst/la0/address_counter[23] , 
        \edb_top_inst/la0/address_counter[24] , \edb_top_inst/la0/address_counter[25] , 
        \edb_top_inst/la0/address_counter[26] , \edb_top_inst/la0/address_counter[27] , 
        \edb_top_inst/la0/opcode[1] , \edb_top_inst/la0/opcode[2] , \edb_top_inst/la0/opcode[3] , 
        \edb_top_inst/la0/bit_count[1] , \edb_top_inst/la0/bit_count[2] , 
        \edb_top_inst/la0/bit_count[3] , \edb_top_inst/la0/bit_count[4] , 
        \edb_top_inst/la0/bit_count[5] , \edb_top_inst/la0/word_count[1] , 
        \edb_top_inst/la0/word_count[2] , \edb_top_inst/la0/word_count[3] , 
        \edb_top_inst/la0/word_count[4] , \edb_top_inst/la0/word_count[5] , 
        \edb_top_inst/la0/word_count[6] , \edb_top_inst/la0/word_count[7] , 
        \edb_top_inst/la0/word_count[8] , \edb_top_inst/la0/word_count[9] , 
        \edb_top_inst/la0/word_count[10] , \edb_top_inst/la0/word_count[11] , 
        \edb_top_inst/la0/word_count[12] , \edb_top_inst/la0/word_count[13] , 
        \edb_top_inst/la0/word_count[14] , \edb_top_inst/la0/word_count[15] , 
        \edb_top_inst/la0/data_out_shift_reg[1] , \edb_top_inst/la0/data_out_shift_reg[2] , 
        \edb_top_inst/la0/data_out_shift_reg[3] , \edb_top_inst/la0/data_out_shift_reg[4] , 
        \edb_top_inst/la0/data_out_shift_reg[5] , \edb_top_inst/la0/data_out_shift_reg[6] , 
        \edb_top_inst/la0/data_out_shift_reg[7] , \edb_top_inst/la0/data_out_shift_reg[8] , 
        \edb_top_inst/la0/data_out_shift_reg[9] , \edb_top_inst/la0/data_out_shift_reg[10] , 
        \edb_top_inst/la0/data_out_shift_reg[11] , \edb_top_inst/la0/data_out_shift_reg[12] , 
        \edb_top_inst/la0/data_out_shift_reg[13] , \edb_top_inst/la0/data_out_shift_reg[14] , 
        \edb_top_inst/la0/data_out_shift_reg[15] , \edb_top_inst/la0/data_out_shift_reg[16] , 
        \edb_top_inst/la0/data_out_shift_reg[17] , \edb_top_inst/la0/data_out_shift_reg[18] , 
        \edb_top_inst/la0/data_out_shift_reg[19] , \edb_top_inst/la0/data_out_shift_reg[20] , 
        \edb_top_inst/la0/data_out_shift_reg[21] , \edb_top_inst/la0/data_out_shift_reg[22] , 
        \edb_top_inst/la0/data_out_shift_reg[23] , \edb_top_inst/la0/data_out_shift_reg[24] , 
        \edb_top_inst/la0/data_out_shift_reg[25] , \edb_top_inst/la0/data_out_shift_reg[26] , 
        \edb_top_inst/la0/data_out_shift_reg[27] , \edb_top_inst/la0/data_out_shift_reg[28] , 
        \edb_top_inst/la0/data_out_shift_reg[29] , \edb_top_inst/la0/data_out_shift_reg[30] , 
        \edb_top_inst/la0/data_out_shift_reg[31] , \edb_top_inst/la0/data_out_shift_reg[32] , 
        \edb_top_inst/la0/data_out_shift_reg[33] , \edb_top_inst/la0/data_out_shift_reg[34] , 
        \edb_top_inst/la0/data_out_shift_reg[35] , \edb_top_inst/la0/data_out_shift_reg[36] , 
        \edb_top_inst/la0/data_out_shift_reg[37] , \edb_top_inst/la0/data_out_shift_reg[38] , 
        \edb_top_inst/la0/data_out_shift_reg[39] , \edb_top_inst/la0/data_out_shift_reg[40] , 
        \edb_top_inst/la0/data_out_shift_reg[41] , \edb_top_inst/la0/data_out_shift_reg[42] , 
        \edb_top_inst/la0/data_out_shift_reg[43] , \edb_top_inst/la0/data_out_shift_reg[44] , 
        \edb_top_inst/la0/data_out_shift_reg[45] , \edb_top_inst/la0/data_out_shift_reg[46] , 
        \edb_top_inst/la0/data_out_shift_reg[47] , \edb_top_inst/la0/data_out_shift_reg[48] , 
        \edb_top_inst/la0/data_out_shift_reg[49] , \edb_top_inst/la0/data_out_shift_reg[50] , 
        \edb_top_inst/la0/data_out_shift_reg[51] , \edb_top_inst/la0/data_out_shift_reg[52] , 
        \edb_top_inst/la0/data_out_shift_reg[53] , \edb_top_inst/la0/data_out_shift_reg[54] , 
        \edb_top_inst/la0/data_out_shift_reg[55] , \edb_top_inst/la0/data_out_shift_reg[56] , 
        \edb_top_inst/la0/data_out_shift_reg[57] , \edb_top_inst/la0/data_out_shift_reg[58] , 
        \edb_top_inst/la0/data_out_shift_reg[59] , \edb_top_inst/la0/data_out_shift_reg[60] , 
        \edb_top_inst/la0/data_out_shift_reg[61] , \edb_top_inst/la0/data_out_shift_reg[62] , 
        \edb_top_inst/la0/data_out_shift_reg[63] , \edb_top_inst/la0/module_state[1] , 
        \edb_top_inst/la0/module_state[2] , \edb_top_inst/la0/module_state[3] , 
        \edb_top_inst/la0/crc_data_out[0] , \edb_top_inst/la0/crc_data_out[1] , 
        \edb_top_inst/la0/crc_data_out[2] , \edb_top_inst/la0/crc_data_out[3] , 
        \edb_top_inst/la0/crc_data_out[4] , \edb_top_inst/la0/crc_data_out[5] , 
        \edb_top_inst/la0/crc_data_out[6] , \edb_top_inst/la0/crc_data_out[7] , 
        \edb_top_inst/la0/crc_data_out[8] , \edb_top_inst/la0/crc_data_out[9] , 
        \edb_top_inst/la0/crc_data_out[10] , \edb_top_inst/la0/crc_data_out[11] , 
        \edb_top_inst/la0/crc_data_out[12] , \edb_top_inst/la0/crc_data_out[13] , 
        \edb_top_inst/la0/crc_data_out[14] , \edb_top_inst/la0/crc_data_out[15] , 
        \edb_top_inst/la0/crc_data_out[16] , \edb_top_inst/la0/crc_data_out[17] , 
        \edb_top_inst/la0/crc_data_out[18] , \edb_top_inst/la0/crc_data_out[19] , 
        \edb_top_inst/la0/crc_data_out[20] , \edb_top_inst/la0/crc_data_out[21] , 
        \edb_top_inst/la0/crc_data_out[22] , \edb_top_inst/la0/crc_data_out[23] , 
        \edb_top_inst/la0/crc_data_out[24] , \edb_top_inst/la0/crc_data_out[25] , 
        \edb_top_inst/la0/crc_data_out[26] , \edb_top_inst/la0/crc_data_out[27] , 
        \edb_top_inst/la0/crc_data_out[28] , \edb_top_inst/la0/crc_data_out[29] , 
        \edb_top_inst/la0/crc_data_out[30] , \edb_top_inst/la0/crc_data_out[31] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/tu_trigger , \edb_top_inst/la0/la_biu_inst/curr_state[0] , 
        \edb_top_inst/la0/la_biu_inst/run_trig_p2 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , \edb_top_inst/la0/la_biu_inst/str_sync , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , \edb_top_inst/la0/la_biu_inst/rdy_sync , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q , \edb_top_inst/la0/data_from_biu[0] , 
        \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] , \edb_top_inst/la0/la_biu_inst/curr_state[3] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[2] , \edb_top_inst/la0/la_biu_inst/curr_state[1] , 
        \edb_top_inst/la0/biu_ready , \edb_top_inst/la0/la_biu_inst/addr_reg[15] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[16] , \edb_top_inst/la0/la_biu_inst/addr_reg[17] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[18] , \edb_top_inst/la0/la_biu_inst/addr_reg[19] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[20] , \edb_top_inst/la0/la_biu_inst/addr_reg[21] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[22] , \edb_top_inst/la0/la_biu_inst/addr_reg[23] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[24] , \edb_top_inst/la0/la_biu_inst/addr_reg[25] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[26] , \edb_top_inst/la0/la_biu_inst/addr_reg[27] , 
        \edb_top_inst/la0/data_from_biu[1] , \edb_top_inst/la0/data_from_biu[2] , 
        \edb_top_inst/la0/data_from_biu[3] , \edb_top_inst/la0/data_from_biu[4] , 
        \edb_top_inst/la0/data_from_biu[5] , \edb_top_inst/la0/data_from_biu[6] , 
        \edb_top_inst/la0/data_from_biu[7] , \edb_top_inst/la0/data_from_biu[8] , 
        \edb_top_inst/la0/data_from_biu[9] , \edb_top_inst/la0/data_from_biu[10] , 
        \edb_top_inst/la0/data_from_biu[11] , \edb_top_inst/la0/data_from_biu[12] , 
        \edb_top_inst/la0/data_from_biu[13] , \edb_top_inst/la0/data_from_biu[14] , 
        \edb_top_inst/la0/data_from_biu[15] , \edb_top_inst/la0/data_from_biu[16] , 
        \edb_top_inst/la0/data_from_biu[17] , \edb_top_inst/la0/data_from_biu[18] , 
        \edb_top_inst/la0/data_from_biu[19] , \edb_top_inst/la0/data_from_biu[20] , 
        \edb_top_inst/la0/data_from_biu[21] , \edb_top_inst/la0/data_from_biu[22] , 
        \edb_top_inst/la0/data_from_biu[23] , \edb_top_inst/la0/data_from_biu[24] , 
        \edb_top_inst/la0/data_from_biu[25] , \edb_top_inst/la0/data_from_biu[26] , 
        \edb_top_inst/la0/data_from_biu[27] , \edb_top_inst/la0/data_from_biu[28] , 
        \edb_top_inst/la0/data_from_biu[29] , \edb_top_inst/la0/data_from_biu[30] , 
        \edb_top_inst/la0/data_from_biu[31] , \edb_top_inst/la0/data_from_biu[32] , 
        \edb_top_inst/la0/data_from_biu[33] , \edb_top_inst/la0/data_from_biu[34] , 
        \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] , 
        \edb_top_inst/la0/la_sample_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 , \edb_top_inst/la0/la_biu_inst/fifo_counter[0] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12] , 
        \edb_top_inst/la0/la_sample_cnt[1] , \edb_top_inst/la0/la_sample_cnt[2] , 
        \edb_top_inst/la0/la_sample_cnt[3] , \edb_top_inst/la0/la_sample_cnt[4] , 
        \edb_top_inst/la0/la_sample_cnt[5] , \edb_top_inst/la0/la_sample_cnt[6] , 
        \edb_top_inst/la0/la_sample_cnt[7] , \edb_top_inst/la0/la_sample_cnt[8] , 
        \edb_top_inst/la0/la_sample_cnt[9] , \edb_top_inst/la0/la_sample_cnt[10] , 
        \edb_top_inst/la0/la_sample_cnt[11] , \edb_top_inst/la0/la_sample_cnt[12] , 
        \edb_top_inst/la0/la_sample_cnt[13] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[1] , \edb_top_inst/la0/la_biu_inst/fifo_counter[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[3] , \edb_top_inst/la0/la_biu_inst/fifo_counter[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[5] , \edb_top_inst/la0/la_biu_inst/fifo_counter[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[7] , \edb_top_inst/la0/la_biu_inst/fifo_counter[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[9] , \edb_top_inst/la0/la_biu_inst/fifo_counter[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[11] , \edb_top_inst/la0/la_biu_inst/fifo_counter[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13] , \edb_top_inst/la0/internal_register_select[1] , 
        \edb_top_inst/la0/internal_register_select[2] , \edb_top_inst/la0/internal_register_select[3] , 
        \edb_top_inst/la0/internal_register_select[4] , \edb_top_inst/la0/internal_register_select[5] , 
        \edb_top_inst/la0/internal_register_select[6] , \edb_top_inst/la0/internal_register_select[7] , 
        \edb_top_inst/la0/internal_register_select[8] , \edb_top_inst/la0/internal_register_select[9] , 
        \edb_top_inst/la0/internal_register_select[10] , \edb_top_inst/la0/internal_register_select[11] , 
        \edb_top_inst/la0/internal_register_select[12] , \edb_top_inst/la0/la_trig_pos[1] , 
        \edb_top_inst/la0/la_trig_pos[2] , \edb_top_inst/la0/la_trig_pos[3] , 
        \edb_top_inst/la0/la_trig_pos[4] , \edb_top_inst/la0/la_trig_pos[5] , 
        \edb_top_inst/la0/la_trig_pos[6] , \edb_top_inst/la0/la_trig_pos[7] , 
        \edb_top_inst/la0/la_trig_pos[8] , \edb_top_inst/la0/la_trig_pos[9] , 
        \edb_top_inst/la0/la_trig_pos[10] , \edb_top_inst/la0/la_trig_pos[11] , 
        \edb_top_inst/la0/la_trig_pos[12] , \edb_top_inst/la0/la_trig_pos[13] , 
        \edb_top_inst/la0/la_trig_pos[14] , \edb_top_inst/la0/la_trig_pos[15] , 
        \edb_top_inst/la0/la_trig_pos[16] , \edb_top_inst/debug_hub_inst/module_id_reg[0] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[1] , \edb_top_inst/debug_hub_inst/module_id_reg[2] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[3] , \edb_top_inst/n60 , 
        \edb_top_inst/n62 , \edb_top_inst/n663 , \edb_top_inst/n665 , 
        \edb_top_inst/n666 , \edb_top_inst/n667 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i6_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i7_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i1_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i2_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i24_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i3_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre , 
        \edb_top_inst/n3117 , \edb_top_inst/n3118 , \edb_top_inst/n3119 , 
        \edb_top_inst/n3120 , \edb_top_inst/n3121 , \edb_top_inst/n3122 , 
        \edb_top_inst/n3123 , \edb_top_inst/n3124 , \edb_top_inst/n3125 , 
        \edb_top_inst/n3126 , \edb_top_inst/n3127 , \edb_top_inst/n3128 , 
        \edb_top_inst/n3129 , \edb_top_inst/n3130 , \edb_top_inst/n3131 , 
        \edb_top_inst/n3132 , \edb_top_inst/n3133 , \edb_top_inst/n3134 , 
        \edb_top_inst/n3135 , \edb_top_inst/n3136 , \edb_top_inst/n3137 , 
        \edb_top_inst/n3138 , \edb_top_inst/n3139 , \edb_top_inst/n3140 , 
        \edb_top_inst/n3141 , \edb_top_inst/n3142 , \edb_top_inst/n3143 , 
        \edb_top_inst/n3144 , \edb_top_inst/n3145 , \edb_top_inst/n3146 , 
        \edb_top_inst/n3147 , \edb_top_inst/n3148 , \edb_top_inst/n3149 , 
        \edb_top_inst/n3150 , \edb_top_inst/n3093 , \edb_top_inst/n3090 , 
        \edb_top_inst/n3151 , \edb_top_inst/n3152 , \edb_top_inst/n3153 , 
        \edb_top_inst/n3154 , \edb_top_inst/n3155 , \edb_top_inst/n3156 , 
        \edb_top_inst/n3157 , \edb_top_inst/n3158 , \edb_top_inst/n3159 , 
        \edb_top_inst/n3160 , \edb_top_inst/n3161 , \edb_top_inst/n3162 , 
        \edb_top_inst/n3163 , \edb_top_inst/n3164 , \edb_top_inst/n3165 , 
        \edb_top_inst/n3166 , \edb_top_inst/n3167 , \edb_top_inst/n3168 , 
        \edb_top_inst/n3169 , \edb_top_inst/n3170 , \edb_top_inst/n3171 , 
        \edb_top_inst/n3172 , \edb_top_inst/n3173 , \edb_top_inst/n3174 , 
        \edb_top_inst/n3175 , \edb_top_inst/n3176 , \edb_top_inst/n3177 , 
        \edb_top_inst/n3178 , \edb_top_inst/n3179 , \edb_top_inst/n3180 , 
        \edb_top_inst/n3181 , \edb_top_inst/n3182 , \edb_top_inst/n3183 , 
        \edb_top_inst/n3184 , \edb_top_inst/n3185 , \edb_top_inst/n3186 , 
        \edb_top_inst/n3187 , \edb_top_inst/n3188 , \edb_top_inst/n3189 , 
        \edb_top_inst/n3190 , \edb_top_inst/n3191 , \edb_top_inst/n3192 , 
        \edb_top_inst/n3193 , \edb_top_inst/n3194 , \edb_top_inst/n3195 , 
        \edb_top_inst/n3196 , \edb_top_inst/n3197 , \edb_top_inst/n3198 , 
        \edb_top_inst/n3199 , \edb_top_inst/n3200 , \edb_top_inst/n1224 , 
        \edb_top_inst/n3201 , \edb_top_inst/n3202 , \edb_top_inst/n3203 , 
        \edb_top_inst/n3204 , \edb_top_inst/n3205 , \edb_top_inst/n3206 , 
        \edb_top_inst/n3207 , \edb_top_inst/n3208 , \edb_top_inst/n3209 , 
        \edb_top_inst/n3210 , \edb_top_inst/n3211 , \edb_top_inst/n3212 , 
        \edb_top_inst/n3213 , \edb_top_inst/n3214 , \edb_top_inst/n3215 , 
        \edb_top_inst/n3216 , \edb_top_inst/n3217 , \edb_top_inst/n3218 , 
        \edb_top_inst/n3219 , \edb_top_inst/n3220 , \edb_top_inst/n3221 , 
        \edb_top_inst/n3222 , \edb_top_inst/n3223 , \edb_top_inst/n3224 , 
        \edb_top_inst/n3225 , \edb_top_inst/n3226 , \edb_top_inst/n3227 , 
        \edb_top_inst/n3228 , \edb_top_inst/n3229 , \edb_top_inst/n3230 , 
        \edb_top_inst/n3231 , \edb_top_inst/n3232 , \edb_top_inst/n3233 , 
        \edb_top_inst/n3234 , \edb_top_inst/n3235 , \edb_top_inst/n3236 , 
        \edb_top_inst/n3237 , \edb_top_inst/n3238 , \edb_top_inst/n3243 , 
        \edb_top_inst/n3244 , \edb_top_inst/n3245 , \edb_top_inst/n3246 , 
        \edb_top_inst/n3247 , \edb_top_inst/n3248 , \edb_top_inst/n3249 , 
        \edb_top_inst/n3250 , \edb_top_inst/n3251 , \edb_top_inst/n3252 , 
        \edb_top_inst/n3253 , \edb_top_inst/n3254 , \edb_top_inst/n3255 , 
        \edb_top_inst/n3256 , \edb_top_inst/n3257 , \edb_top_inst/n3258 , 
        \edb_top_inst/n3259 , \edb_top_inst/n3260 , \edb_top_inst/n3261 , 
        \edb_top_inst/n3262 , \edb_top_inst/n3263 , \edb_top_inst/n3264 , 
        \edb_top_inst/n3265 , \edb_top_inst/n3266 , \edb_top_inst/n3267 , 
        \edb_top_inst/n3268 , \edb_top_inst/n3269 , \edb_top_inst/n3270 , 
        \edb_top_inst/n3271 , \edb_top_inst/n3272 , \edb_top_inst/n3273 , 
        \edb_top_inst/n3274 , \edb_top_inst/n3275 , \edb_top_inst/n3276 , 
        \edb_top_inst/n3277 , \edb_top_inst/n3278 , \edb_top_inst/n3279 , 
        \edb_top_inst/n3280 , \edb_top_inst/n3281 , \edb_top_inst/n3282 , 
        \edb_top_inst/n3283 , \edb_top_inst/n3284 , \edb_top_inst/n3285 , 
        \edb_top_inst/n3286 , \edb_top_inst/n3287 , \edb_top_inst/n3288 , 
        \edb_top_inst/n3289 , \edb_top_inst/n3290 , \edb_top_inst/n3291 , 
        \edb_top_inst/n3292 , \edb_top_inst/n3293 , \edb_top_inst/n3294 , 
        \edb_top_inst/n3295 , \edb_top_inst/n3296 , \edb_top_inst/n3297 , 
        \edb_top_inst/n3298 , \edb_top_inst/n3299 , \edb_top_inst/n3300 , 
        \edb_top_inst/n3301 , \edb_top_inst/n3302 , \edb_top_inst/n3303 , 
        \edb_top_inst/n3304 , \edb_top_inst/n3305 , \edb_top_inst/n3306 , 
        \edb_top_inst/n3307 , \edb_top_inst/n3308 , \edb_top_inst/n3309 , 
        \edb_top_inst/n3310 , \edb_top_inst/n3311 , \edb_top_inst/n3312 , 
        \edb_top_inst/n3313 , \edb_top_inst/n3314 , \edb_top_inst/n3315 , 
        \edb_top_inst/n3316 , \edb_top_inst/n3317 , \edb_top_inst/n3318 , 
        \edb_top_inst/n3319 , \edb_top_inst/n3320 , \edb_top_inst/n3321 , 
        \edb_top_inst/n3322 , \edb_top_inst/n3323 , \edb_top_inst/n3324 , 
        \edb_top_inst/n3325 , \edb_top_inst/n3326 , \edb_top_inst/n3327 , 
        \edb_top_inst/n3328 , \edb_top_inst/n3329 , \edb_top_inst/n3330 , 
        \edb_top_inst/n3331 , \edb_top_inst/n3332 , \edb_top_inst/n3333 , 
        \edb_top_inst/n3334 , \edb_top_inst/n3335 , \edb_top_inst/n3336 , 
        \edb_top_inst/n3337 , \edb_top_inst/n3338 , \edb_top_inst/n3339 , 
        \edb_top_inst/n3340 , \edb_top_inst/n3341 , \edb_top_inst/n3342 , 
        \edb_top_inst/n3343 , \edb_top_inst/n3344 , \edb_top_inst/n3345 , 
        \edb_top_inst/n3346 , \edb_top_inst/n3347 , \edb_top_inst/n3348 , 
        \edb_top_inst/n3349 , \edb_top_inst/n3350 , \edb_top_inst/n3351 , 
        \edb_top_inst/n3352 , \edb_top_inst/n3353 , \edb_top_inst/n3354 , 
        \edb_top_inst/n3355 , \edb_top_inst/n3356 , \edb_top_inst/n3357 , 
        \edb_top_inst/n3358 , \edb_top_inst/n3359 , \edb_top_inst/n3360 , 
        \edb_top_inst/n3361 , \edb_top_inst/n3362 , \edb_top_inst/n3363 , 
        \edb_top_inst/n3364 , \edb_top_inst/n3365 , \edb_top_inst/n3366 , 
        \edb_top_inst/n3367 , \edb_top_inst/n3368 , \edb_top_inst/n3369 , 
        \edb_top_inst/n3370 , \edb_top_inst/n3371 , \edb_top_inst/n3372 , 
        \edb_top_inst/n3373 , \edb_top_inst/n3374 , \edb_top_inst/n3375 , 
        \edb_top_inst/n3376 , \edb_top_inst/n3377 , \edb_top_inst/n3378 , 
        \edb_top_inst/n3379 , \edb_top_inst/n3380 , \edb_top_inst/n3381 , 
        \edb_top_inst/n3382 , \edb_top_inst/n3383 , \edb_top_inst/n3384 , 
        \edb_top_inst/n3385 , \edb_top_inst/n3386 , \edb_top_inst/n3387 , 
        \edb_top_inst/n3388 , \edb_top_inst/n3389 , \edb_top_inst/n3390 , 
        \edb_top_inst/n3391 , \edb_top_inst/n3392 , \edb_top_inst/n3393 , 
        \edb_top_inst/n3394 , \edb_top_inst/n3395 , \edb_top_inst/n3396 , 
        \edb_top_inst/n3397 , \edb_top_inst/n3398 , \edb_top_inst/n3399 , 
        \edb_top_inst/n3400 , \edb_top_inst/n3401 , \edb_top_inst/n3402 , 
        \edb_top_inst/n3403 , \edb_top_inst/n3404 , \edb_top_inst/n3405 , 
        \edb_top_inst/n3406 , \edb_top_inst/n3407 , \edb_top_inst/n3408 , 
        \edb_top_inst/n3409 , \edb_top_inst/n3410 , \edb_top_inst/n3411 , 
        \edb_top_inst/n3412 , \edb_top_inst/n3413 , \edb_top_inst/n3414 , 
        \edb_top_inst/n3415 , \edb_top_inst/n3416 , \edb_top_inst/n3417 , 
        \edb_top_inst/n3418 , \edb_top_inst/n3419 , \edb_top_inst/n3420 , 
        \edb_top_inst/n3421 , \edb_top_inst/n3422 , \edb_top_inst/n3423 , 
        \edb_top_inst/n3424 , \edb_top_inst/n3425 , \edb_top_inst/n3426 , 
        \edb_top_inst/n3427 , \edb_top_inst/n3428 , \edb_top_inst/n3429 , 
        \edb_top_inst/n3430 , \edb_top_inst/n3431 , \edb_top_inst/n3432 , 
        \edb_top_inst/n3433 , \edb_top_inst/n3434 , \edb_top_inst/n3435 , 
        \edb_top_inst/n3436 , \edb_top_inst/n3437 , \edb_top_inst/n3438 , 
        \edb_top_inst/n3439 , \edb_top_inst/n3440 , \edb_top_inst/n3441 , 
        \edb_top_inst/n3442 , \edb_top_inst/n3443 , \edb_top_inst/n3444 , 
        \edb_top_inst/n3445 , \edb_top_inst/n3446 , \edb_top_inst/n3447 , 
        \edb_top_inst/n3448 , \edb_top_inst/n3449 , \edb_top_inst/n3450 , 
        \edb_top_inst/n3451 , \edb_top_inst/n3452 , \edb_top_inst/n3453 , 
        \edb_top_inst/n3454 , \edb_top_inst/n3455 , \edb_top_inst/n3456 , 
        \edb_top_inst/n3457 , \edb_top_inst/n3458 , \edb_top_inst/n3459 , 
        \edb_top_inst/n3460 , \edb_top_inst/n3461 , \edb_top_inst/n3462 , 
        \edb_top_inst/n3463 , \edb_top_inst/n3464 , \edb_top_inst/n3465 , 
        \edb_top_inst/n3466 , \edb_top_inst/n3467 , \edb_top_inst/n3468 , 
        \edb_top_inst/n3469 , \edb_top_inst/n3470 , \edb_top_inst/n3471 , 
        \edb_top_inst/n3472 , \edb_top_inst/n3473 , \edb_top_inst/n3474 , 
        \edb_top_inst/n3475 , \edb_top_inst/n3476 , \edb_top_inst/n3477 , 
        \edb_top_inst/n3478 , \edb_top_inst/n3479 , \edb_top_inst/n3480 , 
        \edb_top_inst/n3481 , \edb_top_inst/n3482 , \edb_top_inst/n3483 , 
        \edb_top_inst/n3484 , \edb_top_inst/n3485 , \edb_top_inst/n3486 , 
        \edb_top_inst/n3487 , \edb_top_inst/n3488 , \edb_top_inst/n3489 , 
        \edb_top_inst/n3490 , \edb_top_inst/n3491 , \edb_top_inst/n3492 , 
        \edb_top_inst/n3493 , \edb_top_inst/n3494 , \edb_top_inst/n3495 , 
        \edb_top_inst/n3496 , \edb_top_inst/n3497 , \edb_top_inst/n3498 , 
        \edb_top_inst/n3499 , \edb_top_inst/n3500 , \edb_top_inst/n3501 , 
        \edb_top_inst/n3502 , \edb_top_inst/n3503 , \edb_top_inst/n3504 , 
        \edb_top_inst/n3505 , \edb_top_inst/n3506 , \edb_top_inst/n3507 , 
        \edb_top_inst/n3508 , \edb_top_inst/n3509 , \edb_top_inst/n3510 , 
        \edb_top_inst/n3511 , \edb_top_inst/n3512 , \edb_top_inst/n3513 , 
        \edb_top_inst/n3514 , \edb_top_inst/n3515 , \edb_top_inst/n3516 , 
        \edb_top_inst/n3517 , \edb_top_inst/n3518 , \edb_top_inst/n3519 , 
        \edb_top_inst/n3520 , \edb_top_inst/n3521 , \edb_top_inst/n3522 , 
        \edb_top_inst/n3523 , \edb_top_inst/n3524 , \edb_top_inst/n3525 , 
        \edb_top_inst/n3526 , \edb_top_inst/n3527 , \edb_top_inst/n3528 , 
        \edb_top_inst/n3529 , \edb_top_inst/n3530 , \edb_top_inst/n3531 , 
        \edb_top_inst/n3532 , \edb_top_inst/n3533 , \edb_top_inst/n3534 , 
        \edb_top_inst/n3535 , \edb_top_inst/n3536 , \edb_top_inst/n3537 , 
        \edb_top_inst/n3538 , \edb_top_inst/n3539 , \edb_top_inst/n3540 , 
        \edb_top_inst/n3541 , \edb_top_inst/n3542 , \edb_top_inst/n3543 , 
        \edb_top_inst/n3544 , \edb_top_inst/n3545 , \edb_top_inst/n3546 , 
        \edb_top_inst/n3547 , \edb_top_inst/n3548 , \edb_top_inst/n3549 , 
        \edb_top_inst/n3550 , \edb_top_inst/n3551 , \edb_top_inst/n3552 , 
        \edb_top_inst/n3553 , \edb_top_inst/n3554 , \edb_top_inst/n3555 , 
        \edb_top_inst/n3556 , \edb_top_inst/n3557 , \edb_top_inst/n3558 , 
        \edb_top_inst/n3559 , \edb_top_inst/n3560 , \edb_top_inst/n3561 , 
        \edb_top_inst/n3562 , \edb_top_inst/n3563 , \edb_top_inst/n3564 , 
        \edb_top_inst/n3565 , \edb_top_inst/n3566 , \edb_top_inst/n3567 , 
        \edb_top_inst/n3568 , \edb_top_inst/n3569 , \edb_top_inst/n3570 , 
        \edb_top_inst/n3571 , \edb_top_inst/n3572 , \edb_top_inst/n3573 , 
        \edb_top_inst/n3574 , \edb_top_inst/n3575 , \edb_top_inst/n3576 , 
        \edb_top_inst/n3577 , \edb_top_inst/n3578 , \edb_top_inst/n3579 , 
        \edb_top_inst/n3580 , \edb_top_inst/n3581 , \edb_top_inst/n3582 , 
        \edb_top_inst/n3583 , \edb_top_inst/n3584 , \edb_top_inst/n3585 , 
        \edb_top_inst/n3586 , \edb_top_inst/n3587 , \edb_top_inst/n3588 , 
        \edb_top_inst/n3589 , \edb_top_inst/n3590 , \edb_top_inst/n3591 , 
        \edb_top_inst/n3592 , \edb_top_inst/n3593 , \edb_top_inst/n3594 , 
        \edb_top_inst/n3595 , \edb_top_inst/n3596 , \edb_top_inst/n3597 , 
        \edb_top_inst/n3598 , \edb_top_inst/n3599 , \edb_top_inst/n3600 , 
        \edb_top_inst/n3601 , \edb_top_inst/n3602 , \edb_top_inst/n3603 , 
        \edb_top_inst/n3604 , \edb_top_inst/n3605 , \edb_top_inst/n3606 , 
        \edb_top_inst/n3607 , \edb_top_inst/n3608 , \edb_top_inst/n3609 , 
        \edb_top_inst/n3610 , \edb_top_inst/n3611 , \edb_top_inst/n3612 , 
        \edb_top_inst/n3613 , \edb_top_inst/n3614 , \edb_top_inst/n3615 , 
        \edb_top_inst/n3616 , \edb_top_inst/n3617 , \edb_top_inst/n3618 , 
        \edb_top_inst/n3619 , \edb_top_inst/n3620 , \edb_top_inst/n3621 , 
        \edb_top_inst/n3622 , \edb_top_inst/n3623 , \edb_top_inst/n3624 , 
        \edb_top_inst/n3625 , \edb_top_inst/n3626 , \edb_top_inst/n3627 , 
        \edb_top_inst/n3628 , \edb_top_inst/n3629 , \edb_top_inst/n3630 , 
        \edb_top_inst/n3631 , \edb_top_inst/n3632 , \edb_top_inst/n3633 , 
        \edb_top_inst/n3634 , \edb_top_inst/n3635 , \edb_top_inst/n3636 , 
        \edb_top_inst/n3637 , \edb_top_inst/n3638 , \edb_top_inst/n3639 , 
        \edb_top_inst/n3640 , \edb_top_inst/n3641 , \edb_top_inst/n3642 , 
        \edb_top_inst/n3643 , \edb_top_inst/n3644 , \edb_top_inst/n3645 , 
        \edb_top_inst/n3646 , \edb_top_inst/n3647 , \edb_top_inst/n3648 , 
        \edb_top_inst/n3649 , \edb_top_inst/n3650 , \edb_top_inst/n3651 , 
        \edb_top_inst/n3652 , \edb_top_inst/n3653 , \edb_top_inst/n3654 , 
        \edb_top_inst/n3655 , \edb_top_inst/n3656 , \edb_top_inst/n3657 , 
        \edb_top_inst/n3658 , \edb_top_inst/n3659 , \edb_top_inst/n3660 , 
        \edb_top_inst/n3661 , \edb_top_inst/n3662 , \edb_top_inst/n3663 , 
        \edb_top_inst/n3664 , \edb_top_inst/n3665 , \edb_top_inst/n3666 , 
        \edb_top_inst/n3667 , \edb_top_inst/n3668 , \edb_top_inst/n3669 , 
        \edb_top_inst/n3670 , \edb_top_inst/n3671 , \edb_top_inst/n3672 , 
        \edb_top_inst/n3673 , \edb_top_inst/n3674 , \edb_top_inst/n3675 , 
        \edb_top_inst/n3676 , \edb_top_inst/n3677 , \edb_top_inst/n3678 , 
        \edb_top_inst/n3679 , \edb_top_inst/n3680 , \edb_top_inst/n3681 , 
        \edb_top_inst/n3682 , \edb_top_inst/n3683 , \edb_top_inst/n3684 , 
        \edb_top_inst/n3685 , \edb_top_inst/n3686 , \edb_top_inst/n3687 , 
        \edb_top_inst/n3688 , \edb_top_inst/n3689 , \edb_top_inst/n3690 , 
        \edb_top_inst/n3691 , \edb_top_inst/n3692 , \edb_top_inst/n3693 , 
        \edb_top_inst/n3694 , \edb_top_inst/n3695 , \edb_top_inst/n3696 , 
        \edb_top_inst/n3697 , \edb_top_inst/n3698 , \edb_top_inst/n3699 , 
        \edb_top_inst/n3096 , n3314, n3315, n3316, n3317, n3318, 
        n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, 
        n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, 
        n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, 
        n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, 
        n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
        n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
        n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, 
        n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, 
        n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, 
        n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, 
        n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
        n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, 
        n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, 
        n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, 
        n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, 
        n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
        n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, 
        n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, 
        n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, 
        n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, 
        n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
        n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, 
        n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
        n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, 
        n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, 
        n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
        n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, 
        n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, 
        n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, 
        n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
        n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
        n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, 
        n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, 
        n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, 
        n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, 
        n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
        n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, 
        n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
        n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, 
        n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, 
        n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, 
        n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, 
        n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, 
        n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, 
        n3671, n3672, n3673, n3689, n3690, n3691, n3692, n3693, 
        n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, 
        n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, 
        n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, 
        n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, 
        n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, 
        n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
        n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, 
        n3750, n3751, n3752, n3753, n3754, wCdcFifoFull, rSRST, 
        \MCsiRxController/MCsi2Decoder/select_39/Select_0/n17 , \MCsiRxController/MCsi2Decoder/n7 , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[0] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qFullAllmost , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE , 
        \MCsiRxController/MCsi2Decoder/n640 , \MCsiRxController/MCsi2Decoder/n659 , 
        \MCsiRxController/MCsi2Decoder/qLineCntRst , \MCsiRxController/MCsi2Decoder/select_39/Select_2/n15 , 
        \MCsiRxController/MCsi2Decoder/select_39/Select_1/n17 , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n21 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n265 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n270 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n275 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n280 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n285 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n290 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n295 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n300 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n305 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n310 , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[1] , \MCsiRxController/MCsi2Decoder/wFtiRd[2] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[3] , \MCsiRxController/MCsi2Decoder/wFtiRd[4] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[5] , \MCsiRxController/MCsi2Decoder/wFtiRd[6] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[7] , \MCsiRxController/MCsi2Decoder/wFtiRd[8] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[9] , \MCsiRxController/MCsi2Decoder/wFtiRd[10] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[11] , \MCsiRxController/MCsi2Decoder/wFtiRd[12] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[13] , \MCsiRxController/MCsi2Decoder/wFtiRd[14] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[15] , \MCsiRxController/MCsi2Decoder/equal_30/n8 , 
        \MCsiRxController/MCsi2Decoder/equal_31/n8 , \MCsiRxController/genblk1[0].mVideoFIFO/qRE , 
        \MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost , \MCsiRxController/genblk1[0].mVideoFIFO/qRVD , 
        \MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 , \MCsiRxController/genblk1[0].mVideoFIFO/n436 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n441 , \MCsiRxController/genblk1[0].mVideoFIFO/n446 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n451 , \MCsiRxController/genblk1[0].mVideoFIFO/n456 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n461 , \MCsiRxController/genblk1[0].mVideoFIFO/n466 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n471 , \MVideoPostProcess/qVtgRstCntCke , 
        \MVideoPostProcess/rVtgRstSel , \MVideoPostProcess/equal_18/n21 , 
        \MVideoPostProcess/inst_adv7511_config/n816 , \MVideoPostProcess/inst_adv7511_config/n833 , 
        \~ceg_net510 , \MVideoPostProcess/inst_adv7511_config/n1107 , \MVideoPostProcess/inst_adv7511_config/n1235 , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] , ceg_net477, 
        ceg_net42, ceg_net1377, \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] , 
        \MVideoPostProcess/inst_adv7511_config/n1243 , \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 , 
        \MVideoPostProcess/rVtgRST[2] , \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 , 
        ceg_net1421, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 , 
        ceg_net1389, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 , 
        ceg_net567, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 , 
        ceg_net1460, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 , 
        ceg_net1523, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 , 
        ceg_net1415, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 , 
        ceg_net617, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] , 
        \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0 , \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 , 
        ceg_net1531, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 , 
        n10449, n10448, n10447, n10446, \MVideoPostProcess/mVideoTimingGen/qVrange , 
        \MVideoPostProcess/inst_adv7511_config/n253 , ceg_net941, \MVideoPostProcess/inst_adv7511_config/n252 , 
        \MVideoPostProcess/inst_adv7511_config/n251 , \MVideoPostProcess/inst_adv7511_config/n250 , 
        \MVideoPostProcess/inst_adv7511_config/n249 , \MVideoPostProcess/inst_adv7511_config/n248 , 
        \MVideoPostProcess/inst_adv7511_config/n247 , \MVideoPostProcess/inst_adv7511_config/n246 , 
        \MVideoPostProcess/inst_adv7511_config/n245 , \MVideoPostProcess/inst_adv7511_config/n244 , 
        \MVideoPostProcess/inst_adv7511_config/n700 , \MVideoPostProcess/inst_adv7511_config/n705 , 
        \MVideoPostProcess/inst_adv7511_config/n710 , \MVideoPostProcess/inst_adv7511_config/n715 , 
        \MVideoPostProcess/inst_adv7511_config/n720 , \MVideoPostProcess/inst_adv7511_config/n725 , 
        \MVideoPostProcess/inst_adv7511_config/n730 , \MVideoPostProcess/inst_adv7511_config/n735 , 
        \MVideoPostProcess/inst_adv7511_config/n740 , \MVideoPostProcess/inst_adv7511_config/n745 , 
        \MVideoPostProcess/inst_adv7511_config/n750 , \MVideoPostProcess/inst_adv7511_config/n755 , 
        \MVideoPostProcess/inst_adv7511_config/n760 , \MVideoPostProcess/inst_adv7511_config/n765 , 
        \MVideoPostProcess/inst_adv7511_config/n770 , \MVideoPostProcess/inst_adv7511_config/n780 , 
        \MVideoPostProcess/inst_adv7511_config/n785 , \MVideoPostProcess/inst_adv7511_config/n790 , 
        \MVideoPostProcess/inst_adv7511_config/n795 , \MVideoPostProcess/inst_adv7511_config/n800 , 
        \MVideoPostProcess/inst_adv7511_config/n805 , \MVideoPostProcess/inst_adv7511_config/n810 , 
        \MVideoPostProcess/mVideoTimingGen/n131 , \MVideoPostProcess/mVideoTimingGen/equal_12/n23 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] , 
        \MVideoPostProcess/mVideoTimingGen/qVde , \MVideoPostProcess/mVideoTimingGen/n267 , 
        \MVideoPostProcess/mVideoTimingGen/rHSync[3] , \MVideoPostProcess/mVideoTimingGen/n130 , 
        \MVideoPostProcess/mVideoTimingGen/n129 , \MVideoPostProcess/mVideoTimingGen/n126 , 
        \MVideoPostProcess/mVideoTimingGen/n125 , \MVideoPostProcess/mVideoTimingGen/n121 , 
        \MVideoPostProcess/mVideoTimingGen/qHrange , \MVideoPostProcess/mVideoTimingGen/rVSync[3] , 
        \MVideoPostProcess/mVideoTimingGen/rVde[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n483 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n488 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n493 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n498 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n503 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n508 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n513 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n518 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n523 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n528 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n533 , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] , 
        \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] , 
        \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] , 
        \genblk1.genblk1[0].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[0].mPulseGenerator/equal_12/n23 , 
        \genblk1.genblk1[1].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[1].mPulseGenerator/n50 , 
        \genblk1.genblk1[3].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[3].mPulseGenerator/n50 , 
        \genblk1.genblk1[4].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[4].mPulseGenerator/n50 , 
        \edb_top_inst/la0/n1325 , \edb_top_inst/ceg_net5 , \edb_top_inst/edb_user_dr[60] , 
        \edb_top_inst/la0/n1297 , \edb_top_inst/la0/n1326 , \edb_top_inst/la0/n1327 , 
        \edb_top_inst/edb_user_dr[62] , \edb_top_inst/edb_user_dr[0] , \edb_top_inst/la0/n1381 , 
        \edb_top_inst/edb_user_dr[42] , \edb_top_inst/la0/n1898 , \edb_top_inst/edb_user_dr[59] , 
        \edb_top_inst/la0/n1950 , \edb_top_inst/la0/data_to_addr_counter[0] , 
        \edb_top_inst/la0/addr_ct_en , \edb_top_inst/edb_user_dr[77] , \edb_top_inst/la0/op_reg_en , 
        \edb_top_inst/la0/n2174 , \edb_top_inst/ceg_net26 , \edb_top_inst/la0/data_to_word_counter[0] , 
        \edb_top_inst/la0/word_ct_en , \edb_top_inst/la0/n2451 , \edb_top_inst/ceg_net14 , 
        \edb_top_inst/la0/module_next_state[0] , \edb_top_inst/la0/n2751 , 
        \edb_top_inst/la0/n3584 , \edb_top_inst/la0/n4417 , \edb_top_inst/la0/n5250 , 
        \edb_top_inst/la0/n6083 , \edb_top_inst/la0/n6972 , \edb_top_inst/la0/n6987 , 
        \edb_top_inst/la0/n7185 , \edb_top_inst/la0/n7869 , \edb_top_inst/la0/n7884 , 
        \edb_top_inst/la0/n8082 , \edb_top_inst/la0/n8710 , \edb_top_inst/la0/n9543 , 
        \edb_top_inst/la0/n10376 , la0_probe10, \edb_top_inst/la0/n11209 , 
        \edb_top_inst/la0/n12042 , \edb_top_inst/la0/n12875 , \edb_top_inst/la0/n13708 , 
        \edb_top_inst/la0/n14541 , \edb_top_inst/la0/n16207 , \edb_top_inst/la0/n17040 , 
        \edb_top_inst/la0/n17887 , \edb_top_inst/la0/n17902 , \edb_top_inst/la0/n18100 , 
        \edb_top_inst/edb_user_dr[64] , \edb_top_inst/la0/regsel_ld_en , 
        \edb_top_inst/edb_user_dr[43] , \edb_top_inst/edb_user_dr[61] , 
        \edb_top_inst/edb_user_dr[63] , \edb_top_inst/edb_user_dr[1] , \edb_top_inst/edb_user_dr[2] , 
        \edb_top_inst/edb_user_dr[3] , \edb_top_inst/edb_user_dr[4] , \edb_top_inst/edb_user_dr[5] , 
        \edb_top_inst/edb_user_dr[6] , \edb_top_inst/edb_user_dr[7] , \edb_top_inst/edb_user_dr[8] , 
        \edb_top_inst/edb_user_dr[9] , \edb_top_inst/edb_user_dr[10] , \edb_top_inst/edb_user_dr[11] , 
        \edb_top_inst/edb_user_dr[12] , \edb_top_inst/edb_user_dr[13] , 
        \edb_top_inst/edb_user_dr[14] , \edb_top_inst/edb_user_dr[15] , 
        \edb_top_inst/edb_user_dr[16] , \edb_top_inst/edb_user_dr[17] , 
        \edb_top_inst/edb_user_dr[18] , \edb_top_inst/edb_user_dr[19] , 
        \edb_top_inst/edb_user_dr[20] , \edb_top_inst/edb_user_dr[21] , 
        \edb_top_inst/edb_user_dr[22] , \edb_top_inst/edb_user_dr[23] , 
        \edb_top_inst/edb_user_dr[24] , \edb_top_inst/edb_user_dr[25] , 
        \edb_top_inst/edb_user_dr[26] , \edb_top_inst/edb_user_dr[27] , 
        \edb_top_inst/edb_user_dr[28] , \edb_top_inst/edb_user_dr[29] , 
        \edb_top_inst/edb_user_dr[30] , \edb_top_inst/edb_user_dr[31] , 
        \edb_top_inst/edb_user_dr[32] , \edb_top_inst/edb_user_dr[33] , 
        \edb_top_inst/edb_user_dr[34] , \edb_top_inst/edb_user_dr[35] , 
        \edb_top_inst/edb_user_dr[36] , \edb_top_inst/edb_user_dr[37] , 
        \edb_top_inst/edb_user_dr[38] , \edb_top_inst/edb_user_dr[39] , 
        \edb_top_inst/edb_user_dr[40] , \edb_top_inst/edb_user_dr[41] , 
        \edb_top_inst/edb_user_dr[44] , \edb_top_inst/edb_user_dr[45] , 
        \edb_top_inst/edb_user_dr[46] , \edb_top_inst/edb_user_dr[47] , 
        \edb_top_inst/edb_user_dr[48] , \edb_top_inst/edb_user_dr[49] , 
        \edb_top_inst/edb_user_dr[50] , \edb_top_inst/edb_user_dr[51] , 
        \edb_top_inst/edb_user_dr[52] , \edb_top_inst/edb_user_dr[53] , 
        \edb_top_inst/edb_user_dr[54] , \edb_top_inst/edb_user_dr[55] , 
        \edb_top_inst/edb_user_dr[56] , \edb_top_inst/edb_user_dr[57] , 
        \edb_top_inst/edb_user_dr[58] , \edb_top_inst/la0/data_to_addr_counter[1] , 
        \edb_top_inst/la0/data_to_addr_counter[2] , \edb_top_inst/la0/data_to_addr_counter[3] , 
        \edb_top_inst/la0/data_to_addr_counter[4] , \edb_top_inst/la0/data_to_addr_counter[5] , 
        \edb_top_inst/la0/data_to_addr_counter[6] , \edb_top_inst/la0/data_to_addr_counter[7] , 
        \edb_top_inst/la0/data_to_addr_counter[8] , \edb_top_inst/la0/data_to_addr_counter[9] , 
        \edb_top_inst/la0/data_to_addr_counter[10] , \edb_top_inst/la0/data_to_addr_counter[11] , 
        \edb_top_inst/la0/data_to_addr_counter[12] , \edb_top_inst/la0/data_to_addr_counter[13] , 
        \edb_top_inst/la0/data_to_addr_counter[14] , \edb_top_inst/la0/data_to_addr_counter[15] , 
        \edb_top_inst/la0/data_to_addr_counter[16] , \edb_top_inst/la0/data_to_addr_counter[17] , 
        \edb_top_inst/la0/data_to_addr_counter[18] , \edb_top_inst/la0/data_to_addr_counter[19] , 
        \edb_top_inst/la0/data_to_addr_counter[20] , \edb_top_inst/la0/data_to_addr_counter[21] , 
        \edb_top_inst/la0/data_to_addr_counter[22] , \edb_top_inst/la0/data_to_addr_counter[23] , 
        \edb_top_inst/la0/data_to_addr_counter[24] , \edb_top_inst/la0/data_to_addr_counter[25] , 
        \edb_top_inst/la0/data_to_addr_counter[26] , \edb_top_inst/la0/data_to_addr_counter[27] , 
        \edb_top_inst/edb_user_dr[78] , \edb_top_inst/edb_user_dr[79] , 
        \edb_top_inst/edb_user_dr[80] , \edb_top_inst/la0/n2173 , \edb_top_inst/la0/n2172 , 
        \edb_top_inst/la0/n2171 , \edb_top_inst/la0/n2170 , \edb_top_inst/la0/n2169 , 
        \edb_top_inst/la0/data_to_word_counter[1] , \edb_top_inst/la0/data_to_word_counter[2] , 
        \edb_top_inst/la0/data_to_word_counter[3] , \edb_top_inst/la0/data_to_word_counter[4] , 
        \edb_top_inst/la0/data_to_word_counter[5] , \edb_top_inst/la0/data_to_word_counter[6] , 
        \edb_top_inst/la0/data_to_word_counter[7] , \edb_top_inst/la0/data_to_word_counter[8] , 
        \edb_top_inst/la0/data_to_word_counter[9] , \edb_top_inst/la0/data_to_word_counter[10] , 
        \edb_top_inst/la0/data_to_word_counter[11] , \edb_top_inst/la0/data_to_word_counter[12] , 
        \edb_top_inst/la0/data_to_word_counter[13] , \edb_top_inst/la0/data_to_word_counter[14] , 
        \edb_top_inst/la0/data_to_word_counter[15] , \edb_top_inst/la0/n2450 , 
        \edb_top_inst/la0/n2449 , \edb_top_inst/la0/n2448 , \edb_top_inst/la0/n2447 , 
        \edb_top_inst/la0/n2446 , \edb_top_inst/la0/n2445 , \edb_top_inst/la0/n2444 , 
        \edb_top_inst/la0/n2443 , \edb_top_inst/la0/n2442 , \edb_top_inst/la0/n2441 , 
        \edb_top_inst/la0/n2440 , \edb_top_inst/la0/n2439 , \edb_top_inst/la0/n2438 , 
        \edb_top_inst/la0/n2437 , \edb_top_inst/la0/n2436 , \edb_top_inst/la0/n2435 , 
        \edb_top_inst/la0/n2434 , \edb_top_inst/la0/n2433 , \edb_top_inst/la0/n2432 , 
        \edb_top_inst/la0/n2431 , \edb_top_inst/la0/n2430 , \edb_top_inst/la0/n2429 , 
        \edb_top_inst/la0/n2428 , \edb_top_inst/la0/n2427 , \edb_top_inst/la0/n2426 , 
        \edb_top_inst/la0/n2425 , \edb_top_inst/la0/n2424 , \edb_top_inst/la0/n2423 , 
        \edb_top_inst/la0/n2422 , \edb_top_inst/la0/n2421 , \edb_top_inst/la0/n2420 , 
        \edb_top_inst/la0/n2419 , \edb_top_inst/la0/n2418 , \edb_top_inst/la0/n2417 , 
        \edb_top_inst/la0/n2416 , \edb_top_inst/la0/n2415 , \edb_top_inst/la0/n2414 , 
        \edb_top_inst/la0/n2413 , \edb_top_inst/la0/n2412 , \edb_top_inst/la0/n2411 , 
        \edb_top_inst/la0/n2410 , \edb_top_inst/la0/n2409 , \edb_top_inst/la0/n2408 , 
        \edb_top_inst/la0/n2407 , \edb_top_inst/la0/n2406 , \edb_top_inst/la0/n2405 , 
        \edb_top_inst/la0/n2404 , \edb_top_inst/la0/n2403 , \edb_top_inst/la0/n2402 , 
        \edb_top_inst/la0/n2401 , \edb_top_inst/la0/n2400 , \edb_top_inst/la0/n2399 , 
        \edb_top_inst/la0/n2398 , \edb_top_inst/la0/n2397 , \edb_top_inst/la0/n2396 , 
        \edb_top_inst/la0/n2395 , \edb_top_inst/la0/n2394 , \edb_top_inst/la0/n2393 , 
        \edb_top_inst/la0/n2392 , \edb_top_inst/la0/n2391 , \edb_top_inst/la0/n2390 , 
        \edb_top_inst/la0/n2389 , \edb_top_inst/la0/n2388 , \edb_top_inst/la0/module_next_state[1] , 
        \edb_top_inst/la0/module_next_state[2] , \edb_top_inst/la0/module_next_state[3] , 
        \edb_top_inst/la0/axi_crc_i/n150 , \edb_top_inst/ceg_net221 , \edb_top_inst/la0/axi_crc_i/n149 , 
        \edb_top_inst/la0/axi_crc_i/n148 , \edb_top_inst/la0/axi_crc_i/n147 , 
        \edb_top_inst/la0/axi_crc_i/n146 , \edb_top_inst/la0/axi_crc_i/n145 , 
        \edb_top_inst/la0/axi_crc_i/n144 , \edb_top_inst/la0/axi_crc_i/n143 , 
        \edb_top_inst/la0/axi_crc_i/n142 , \edb_top_inst/la0/axi_crc_i/n141 , 
        \edb_top_inst/la0/axi_crc_i/n140 , \edb_top_inst/la0/axi_crc_i/n139 , 
        \edb_top_inst/la0/axi_crc_i/n138 , \edb_top_inst/la0/axi_crc_i/n137 , 
        \edb_top_inst/la0/axi_crc_i/n136 , \edb_top_inst/la0/axi_crc_i/n135 , 
        \edb_top_inst/la0/axi_crc_i/n134 , \edb_top_inst/la0/axi_crc_i/n133 , 
        \edb_top_inst/la0/axi_crc_i/n132 , \edb_top_inst/la0/axi_crc_i/n131 , 
        \edb_top_inst/la0/axi_crc_i/n130 , \edb_top_inst/la0/axi_crc_i/n129 , 
        \edb_top_inst/la0/axi_crc_i/n128 , \edb_top_inst/la0/axi_crc_i/n127 , 
        \edb_top_inst/la0/axi_crc_i/n126 , \edb_top_inst/la0/axi_crc_i/n125 , 
        \edb_top_inst/la0/axi_crc_i/n124 , \edb_top_inst/la0/axi_crc_i/n123 , 
        \edb_top_inst/la0/axi_crc_i/n122 , \edb_top_inst/la0/axi_crc_i/n121 , 
        \edb_top_inst/la0/axi_crc_i/n120 , \edb_top_inst/la0/axi_crc_i/n119 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n41 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n50 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n38 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n36 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n34 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n21 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n15 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n41 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n50 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n21 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n15 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n15374 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n10 , \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n17 , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/equal_9/n3 , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n26 , \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n15 , 
        \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n9 , \edb_top_inst/la0/trigger_tu/n131 , 
        \edb_top_inst/la0/la_biu_inst/next_state[0] , \edb_top_inst/la0/la_biu_inst/run_trig_p1 , 
        \edb_top_inst/la0/la_biu_inst/n374 , \edb_top_inst/la0/la_biu_inst/n1303 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[0] , \edb_top_inst/la0/la_biu_inst/next_fsm_state[0] , 
        \edb_top_inst/ceg_net351 , \edb_top_inst/la0/la_biu_inst/n1288 , 
        \edb_top_inst/la0/n25424 , \edb_top_inst/la0/la_biu_inst/next_state[2] , 
        \edb_top_inst/la0/la_biu_inst/next_state[1] , \edb_top_inst/ceg_net348 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[3] , \edb_top_inst/la0/la_biu_inst/fifo_dout[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[5] , \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[7] , \edb_top_inst/la0/la_biu_inst/fifo_dout[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[9] , \edb_top_inst/la0/la_biu_inst/fifo_dout[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[11] , \edb_top_inst/la0/la_biu_inst/fifo_dout[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[13] , \edb_top_inst/la0/la_biu_inst/fifo_dout[14] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[15] , \edb_top_inst/la0/la_biu_inst/fifo_dout[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[17] , \edb_top_inst/la0/la_biu_inst/fifo_dout[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[19] , \edb_top_inst/la0/la_biu_inst/fifo_dout[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[21] , \edb_top_inst/la0/la_biu_inst/fifo_dout[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[23] , \edb_top_inst/la0/la_biu_inst/fifo_dout[24] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[25] , \edb_top_inst/la0/la_biu_inst/fifo_dout[26] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[27] , \edb_top_inst/la0/la_biu_inst/fifo_dout[28] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[29] , \edb_top_inst/la0/la_biu_inst/fifo_dout[30] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[31] , \edb_top_inst/la0/la_biu_inst/fifo_dout[32] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[33] , \edb_top_inst/la0/la_biu_inst/fifo_dout[34] , 
        \edb_top_inst/la0/la_biu_inst/next_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , 
        \edb_top_inst/la0/la_biu_inst/fifo_rstn , \edb_top_inst/la0/la_biu_inst/n2043 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 , \edb_top_inst/la0/la_biu_inst/fifo_push , 
        \edb_top_inst/ceg_net355 , \edb_top_inst/n1019 , \edb_top_inst/n1017 , 
        \edb_top_inst/n1015 , \edb_top_inst/n1013 , \edb_top_inst/n1011 , 
        \edb_top_inst/n1009 , \edb_top_inst/n1007 , \edb_top_inst/n1005 , 
        \edb_top_inst/n1003 , \edb_top_inst/n1001 , \edb_top_inst/n999 , 
        \edb_top_inst/n998 , \edb_top_inst/n662 , \edb_top_inst/n996 , 
        \edb_top_inst/n994 , \edb_top_inst/n992 , \edb_top_inst/n990 , 
        \edb_top_inst/n988 , \edb_top_inst/n986 , \edb_top_inst/n984 , 
        \edb_top_inst/n981 , \edb_top_inst/n978 , \edb_top_inst/n976 , 
        \edb_top_inst/n974 , \edb_top_inst/n664 , \edb_top_inst/n971 , 
        \edb_top_inst/n969 , \edb_top_inst/n967 , \edb_top_inst/n965 , 
        \edb_top_inst/n963 , \edb_top_inst/n961 , \edb_top_inst/n959 , 
        \edb_top_inst/n957 , \edb_top_inst/n955 , \edb_top_inst/n953 , 
        \edb_top_inst/n951 , \edb_top_inst/n877 , \edb_top_inst/n900 , 
        \edb_top_inst/n898 , \edb_top_inst/n896 , \edb_top_inst/n894 , 
        \edb_top_inst/n892 , \edb_top_inst/n890 , \edb_top_inst/n888 , 
        \edb_top_inst/n886 , \edb_top_inst/n884 , \edb_top_inst/n882 , 
        \edb_top_inst/n880 , \edb_top_inst/n879 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[12] , 
        \edb_top_inst/n878 , \edb_top_inst/n923 , \edb_top_inst/n921 , 
        \edb_top_inst/n919 , \edb_top_inst/n917 , \edb_top_inst/n915 , 
        \edb_top_inst/n913 , \edb_top_inst/n911 , \edb_top_inst/n909 , 
        \edb_top_inst/n907 , \edb_top_inst/n905 , \edb_top_inst/n903 , 
        \edb_top_inst/n902 , \edb_top_inst/edb_user_dr[65] , \edb_top_inst/edb_user_dr[66] , 
        \edb_top_inst/edb_user_dr[67] , \edb_top_inst/edb_user_dr[68] , 
        \edb_top_inst/edb_user_dr[69] , \edb_top_inst/edb_user_dr[70] , 
        \edb_top_inst/edb_user_dr[71] , \edb_top_inst/edb_user_dr[72] , 
        \edb_top_inst/edb_user_dr[73] , \edb_top_inst/edb_user_dr[74] , 
        \edb_top_inst/edb_user_dr[75] , \edb_top_inst/edb_user_dr[76] , 
        \edb_top_inst/debug_hub_inst/n266 , \edb_top_inst/debug_hub_inst/n95 , 
        \edb_top_inst/edb_user_dr[81] , \edb_top_inst/n881 , \edb_top_inst/n883 , 
        \edb_top_inst/n885 , \edb_top_inst/n887 , \edb_top_inst/n889 , 
        \edb_top_inst/n891 , \edb_top_inst/n893 , \edb_top_inst/n895 , 
        \edb_top_inst/n897 , \edb_top_inst/n899 , \edb_top_inst/n901 , 
        \edb_top_inst/n904 , \edb_top_inst/n906 , \edb_top_inst/n908 , 
        \edb_top_inst/n910 , \edb_top_inst/n912 , \edb_top_inst/n914 , 
        \edb_top_inst/n916 , \edb_top_inst/n918 , \edb_top_inst/n920 , 
        \edb_top_inst/n922 , \edb_top_inst/n924 , \edb_top_inst/n954 , 
        \edb_top_inst/n956 , \edb_top_inst/n958 , \edb_top_inst/n960 , 
        \edb_top_inst/n962 , \edb_top_inst/n964 , \edb_top_inst/n966 , 
        \edb_top_inst/n968 , \edb_top_inst/n970 , \edb_top_inst/n972 , 
        \edb_top_inst/n977 , \edb_top_inst/n979 , \edb_top_inst/n982 , 
        \edb_top_inst/n985 , \edb_top_inst/n987 , \edb_top_inst/n989 , 
        \edb_top_inst/n991 , \edb_top_inst/n993 , \edb_top_inst/n995 , 
        \edb_top_inst/n997 , \edb_top_inst/n1000 , \edb_top_inst/n1002 , 
        \edb_top_inst/n1004 , \edb_top_inst/n1006 , \edb_top_inst/n1008 , 
        \edb_top_inst/n1010 , \edb_top_inst/n1012 , \edb_top_inst/n1014 , 
        \edb_top_inst/n1016 , \edb_top_inst/n1018 , \edb_top_inst/n1020 , 
        \edb_top_inst/n1023 , \edb_top_inst/n1025 , \edb_top_inst/n1027 , 
        \edb_top_inst/n1038 , \edb_top_inst/n1040 , \edb_top_inst/n1042 , 
        \edb_top_inst/n1044 , \edb_top_inst/n1046 , \edb_top_inst/n1048 , 
        \edb_top_inst/n1050 , \edb_top_inst/n1052 , \edb_top_inst/n1054 , 
        \edb_top_inst/n1056 , \edb_top_inst/n1058 , \edb_top_inst/n1060 , 
        \edb_top_inst/n1062 , \edb_top_inst/n1064 , \edb_top_inst/n1066 , 
        \edb_top_inst/n1068 , \edb_top_inst/n1070 , \edb_top_inst/n1072 , 
        \edb_top_inst/n1074 , \edb_top_inst/n1076 , \edb_top_inst/n1078 , 
        \edb_top_inst/n1080 , \edb_top_inst/n1082 , \edb_top_inst/n1084 , 
        \edb_top_inst/n1086 , \edb_top_inst/n1088 , \edb_top_inst/n1099 , 
        \edb_top_inst/n1101 , \edb_top_inst/n1103 , \edb_top_inst/n1105 , 
        \edb_top_inst/n1107 , \edb_top_inst/n1109 , \edb_top_inst/n1111 , 
        \edb_top_inst/n1116 , \edb_top_inst/n1118 , \edb_top_inst/n1120 , 
        \edb_top_inst/n1203 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , \edb_top_inst/n3115 , 
        \edb_top_inst/n59 , \edb_top_inst/n1087 , \edb_top_inst/n1085 , 
        \edb_top_inst/n1083 , \edb_top_inst/n1081 , \edb_top_inst/n1079 , 
        \edb_top_inst/n1077 , \edb_top_inst/n1075 , \edb_top_inst/n1073 , 
        \edb_top_inst/n1071 , \edb_top_inst/n1069 , \edb_top_inst/n1067 , 
        \edb_top_inst/n1065 , \edb_top_inst/n1063 , \edb_top_inst/n1061 , 
        \edb_top_inst/n1059 , \edb_top_inst/n1057 , \edb_top_inst/n1202 , 
        \edb_top_inst/n1055 , \edb_top_inst/n1119 , \edb_top_inst/n1053 , 
        \edb_top_inst/n1117 , \edb_top_inst/n1051 , \edb_top_inst/n1115 , 
        \edb_top_inst/n1049 , \edb_top_inst/n1110 , \edb_top_inst/n1047 , 
        \edb_top_inst/n1108 , \edb_top_inst/n1045 , \edb_top_inst/n1106 , 
        \edb_top_inst/n1043 , \edb_top_inst/n1104 , \edb_top_inst/n1041 , 
        \edb_top_inst/n1102 , \edb_top_inst/n1039 , \edb_top_inst/n1100 , 
        \edb_top_inst/n1037 , \edb_top_inst/n1098 , \edb_top_inst/n1035 , 
        \edb_top_inst/n1096 , \edb_top_inst/n61 , \edb_top_inst/n1026 , 
        \edb_top_inst/n1024 , \edb_top_inst/n1022 , \edb_top_inst/n1021 , 
        n9781, n9980, n10054, n10055, n10056, n10057, n10058, 
        n10059, n10060, n10061, n10062, n10063, n10064, n10065, 
        n10066, n10067, n10068, n10069, n10070, n10071, n10072, 
        n10073, n10074, n10075, n10076, n10077, n10078, n10079, 
        n10080, n10081, n10082, n10083, n10084, n10085, n10086, 
        n10087, n10088, n10089, n10090, n10091, n10092, n10093, 
        n10094, n10095, n10096, n10097, n10098, n10099, n10100, 
        n10101, n10102, n10103, n10104, n10105, n10106, n10107, 
        n10108, n10109, n10110, n10111, n10112, n10113, n10114, 
        n10115, n10116, n10117, n10118, n10119, n10120, n10121, 
        n10122, n10123, n10124, n10126, n10127, n10128, n10129, 
        n10130, n10131, n10132, n10133, n10134, n10135, n10136, 
        n10137, n10138, n10139, n10140, n10141, n10142, n10143, 
        n10144, n10145, n10146, n10147, n10148, n10149, n10150, 
        n10151, n10152, n10153, n10154, n10155, n10156, n10157, 
        n10158, n10159, n10160, n10161, n10162, n10163, n10164, 
        n10165, n10166, n10167, n10168, n10169, n10170, n10171, 
        n10172, n10173, n10174, n10175, n10176, n10177, n10178, 
        n10179, n10180, n10181, n10182, n10183, n10184, n10185, 
        n10186, n10187, n10188, n10189, n10190, n10191, n10192, 
        n10193, n10194, n10195, n10196, n10197, n10198, n10199, 
        n10201, n10203, n10204, n10205, n10206, n10207, n10208, 
        n10209, n10210, n10211, n10212, n10213, n10214, n10220, 
        n10221, n10222, n10223, n10224, n10225, n10226, n10227, 
        n10228, n10229, n10230, n10231, n10232, n10233, n10234, 
        n10235, n10236, n10237, n10238, n10239, n10240, n10241, 
        n10242, n10243, n10244, n10245, n10246, n10247, n10248, 
        n10249, n10250, n10251, n10252, n10253, n10254, n10255, 
        n10256, n10257, n10258, n10259, n10260, n10261, n10262, 
        n10263, n10264, n10265, n10266, n10267, n10268, n10269, 
        n10270, n10271, n10272, n10273, n10274, n10275, n10276, 
        n10277, n10278, n10279, n10280, n10281, n10282, n10283, 
        n10284, n10285, n10286, n10287, n10288, n10289, n10290, 
        n10291, n10292, n10293, n10294, n10295, n10296, n10297, 
        n10298, n10299, n10300, n10301, n10302, n10303, n10304, 
        n10305, n10306, n10307, n10308, n10309, n10310, n10311, 
        n10312, n10313, n10314, n10315, n10316, n10317, n10318, 
        n10319, n10320, n10321, n10322, n10323, n10324, n10325, 
        n10326, n10327, n10328, n10329, n10330, n10331, n10332, 
        n10333, n10334, n10335, n10336, n10337, n10338, n10339, 
        n10340, n10341, n10342, n10343, n10344, n10345, n10346, 
        n10347, n10348, n10349, n10350, n10351, n10352, n10353, 
        n10354, n10355, n10356, n10357, n10358, n10359, n10360, 
        n10361, n10362, n10363, n10364, n10365, n10366, n10367, 
        n10368, n10369, n10370, n10371, n10372, n10373, n10374, 
        n10375, n10376, n10377, n10378, n10379, n10380, n10381, 
        n10382, n10383, n10384, n10385, n10386, n10387, n10388, 
        n10389, n10390, n10391, n10392, n10393, n10394, n10395, 
        n10396, n10397, n10398, n10399, n10400, n10401, n10402, 
        n10403, n10404, n10405, n10406, n10407, n10408, n10409, 
        n10410, n10411, n10412, n10413, n10414, n10415, n10416, 
        n10417, n10418, n10419, n10420, n10421, n10422, n10423, 
        n10424, n10425, n10426, n10427, n10428, n10429, n10430, 
        n10431, n10432, n10433, n10434, n10435, n10436, n10437, 
        n10438, n10439, n10440, n10441, n10442, n10443, n10444, 
        n10445;
    
    assign MipiDphyRx1_RST0_N = MipiDphyRx1_RESET_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[2] = MipiDphyRx1_STOPSTATE_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_REQUEST_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TURN_REQUEST = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_FORCE_RX_MODE = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[7] = MipiDphyRx1_RX_CLK_ACTIVE_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[10] = MipiDphyRx1_RX_ACTIVE_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[24] = MipiDphyRx1_RX_VALID_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[25] = MipiDphyRx1_RX_VALID_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[0] = MipiDphyRx1_RX_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[3] = MipiDphyRx1_RX_SKEW_CAL_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[4] = MipiDphyRx1_RX_DATA_HS_LAN0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_LPDT_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_VALID_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_ULPS_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[17] = MipiDphyRx1_WORD_CLKOUT_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[1] = MipiDphyRx1_RX_CLK_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_CLK_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign pll_inst1_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[23] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[22] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[21] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[20] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[19] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[18] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[16] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[15] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[14] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[13] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[12] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[11] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[9] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[8] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign jtag_inst1_TDO = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign pll_inst2_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_CELL_NAME=VCC */ ;
    assign MipiDphyRx1_TX_ULPS_EXIT = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_FF \MipiDphyRx1_RST0_N~FF  (.D(oLed[0]), .CE(1'b1), .CLK(iSCLK), 
           .SR(iPushSw[0]), .Q(MipiDphyRx1_RESET_N)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MTopTi180MIPI25GRxHDMIV101.v(142)
    defparam \MipiDphyRx1_RST0_N~FF .CLK_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RST0_N~FF .CE_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RST0_N~FF .SR_POLARITY = 1'b0;
    defparam \MipiDphyRx1_RST0_N~FF .D_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RST0_N~FF .SR_SYNC = 1'b0;
    defparam \MipiDphyRx1_RST0_N~FF .SR_VALUE = 1'b0;
    defparam \MipiDphyRx1_RST0_N~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rBRST~FF  (.D(oLed[0]), .CE(1'b1), .CLK(iBCLK), .SR(iPushSw[0]), 
           .Q(rBRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MTopTi180MIPI25GRxHDMIV101.v(149)
    defparam \rBRST~FF .CLK_POLARITY = 1'b1;
    defparam \rBRST~FF .CE_POLARITY = 1'b1;
    defparam \rBRST~FF .SR_POLARITY = 1'b0;
    defparam \rBRST~FF .D_POLARITY = 1'b0;
    defparam \rBRST~FF .SR_SYNC = 1'b0;
    defparam \rBRST~FF .SR_VALUE = 1'b1;
    defparam \rBRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rVRST~FF  (.D(oLed[0]), .CE(1'b1), .CLK(iVCLK), .SR(iPushSw[0]), 
           .Q(rVRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MTopTi180MIPI25GRxHDMIV101.v(160)
    defparam \rVRST~FF .CLK_POLARITY = 1'b1;
    defparam \rVRST~FF .CE_POLARITY = 1'b1;
    defparam \rVRST~FF .SR_POLARITY = 1'b0;
    defparam \rVRST~FF .D_POLARITY = 1'b0;
    defparam \rVRST~FF .SR_SYNC = 1'b0;
    defparam \rVRST~FF .SR_VALUE = 1'b1;
    defparam \rVRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rnVRST~FF  (.D(oLed[0]), .CE(1'b1), .CLK(iVCLK), .SR(iPushSw[0]), 
           .Q(rnVRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MTopTi180MIPI25GRxHDMIV101.v(164)
    defparam \rnVRST~FF .CLK_POLARITY = 1'b1;
    defparam \rnVRST~FF .CE_POLARITY = 1'b1;
    defparam \rnVRST~FF .SR_POLARITY = 1'b0;
    defparam \rnVRST~FF .D_POLARITY = 1'b1;
    defparam \rnVRST~FF .SR_SYNC = 1'b0;
    defparam \rnVRST~FF .SR_VALUE = 1'b0;
    defparam \rnVRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[3]~FF  (.D(1'b1), .CE(wCdcFifoFull), .CLK(iSCLK), .SR(rSRST), 
           .Q(oLed[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MTopTi180MIPI25GRxHDMIV101.v(368)
    defparam \oLed[3]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[3]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[3]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[3]~FF .D_POLARITY = 1'b1;
    defparam \oLed[3]~FF .SR_SYNC = 1'b1;
    defparam \oLed[3]~FF .SR_VALUE = 1'b0;
    defparam \oLed[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe18[0]~FF  (.D(oTestPort[0]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\la0_probe18[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe18[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe18[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe18[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe18[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe18[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe18[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe18[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/select_39/Select_0/n17 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\MCsiRxController/MCsi2Decoder/rHsSt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(226)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs~FF  (.D(MipiDphyRx1_RX_SYNC_HS_LAN1), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF  (.D(\MCsiRxController/MCsi2Decoder/n7 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rSRST_2~FF  (.D(oLed[0]), .CE(1'b1), .CLK(iSCLK), .SR(iPushSw[0]), 
           .Q(rSRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MTopTi180MIPI25GRxHDMIV101.v(138)
    defparam \rSRST_2~FF .CLK_POLARITY = 1'b1;
    defparam \rSRST_2~FF .CE_POLARITY = 1'b1;
    defparam \rSRST_2~FF .SR_POLARITY = 1'b0;
    defparam \rSRST_2~FF .D_POLARITY = 1'b0;
    defparam \rSRST_2~FF .SR_SYNC = 1'b0;
    defparam \rSRST_2~FF .SR_VALUE = 1'b1;
    defparam \rSRST_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe15~FF  (.D(MipiDphyRx1_STOPSTATE_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(la0_probe15)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe15~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe15~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe15~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe15~FF .D_POLARITY = 1'b1;
    defparam \la0_probe15~FF .SR_SYNC = 1'b0;
    defparam \la0_probe15~FF .SR_VALUE = 1'b0;
    defparam \la0_probe15~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe2~FF  (.D(MipiDphyRx1_ERR_ESC_LAN0), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(la0_probe2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe2~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe2~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe2~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe2~FF .D_POLARITY = 1'b1;
    defparam \la0_probe2~FF .SR_SYNC = 1'b0;
    defparam \la0_probe2~FF .SR_VALUE = 1'b0;
    defparam \la0_probe2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe0~FF  (.D(MipiDphyRx1_ERR_CONTROL_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(la0_probe0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe0~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe0~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe0~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe0~FF .D_POLARITY = 1'b1;
    defparam \la0_probe0~FF .SR_SYNC = 1'b0;
    defparam \la0_probe0~FF .SR_VALUE = 1'b0;
    defparam \la0_probe0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe16~FF  (.D(MipiDphyRx1_RX_TRIGGER_ESC[0]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(la0_probe16)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe16~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe16~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe16~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe16~FF .D_POLARITY = 1'b1;
    defparam \la0_probe16~FF .SR_SYNC = 1'b0;
    defparam \la0_probe16~FF .SR_VALUE = 1'b0;
    defparam \la0_probe16~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe4~FF  (.D(MipiDphyRx1_DIRECTION), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(la0_probe4)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe4~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe4~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe4~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe4~FF .D_POLARITY = 1'b1;
    defparam \la0_probe4~FF .SR_SYNC = 1'b0;
    defparam \la0_probe4~FF .SR_VALUE = 1'b0;
    defparam \la0_probe4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe1~FF  (.D(MipiDphyRx1_ERR_CONTENTION_LP0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(la0_probe1)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe1~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe1~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe1~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe1~FF .D_POLARITY = 1'b1;
    defparam \la0_probe1~FF .SR_SYNC = 1'b0;
    defparam \la0_probe1~FF .SR_VALUE = 1'b0;
    defparam \la0_probe1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8~FF  (.D(MipiDphyRx1_ERR_CONTENTION_LP1), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(la0_probe8)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe8~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe12~FF  (.D(la0_probe12), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(la0_probe12)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe12~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe12~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe12~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe12~FF .D_POLARITY = 1'b0;
    defparam \la0_probe12~FF .SR_SYNC = 1'b0;
    defparam \la0_probe12~FF .SR_VALUE = 1'b0;
    defparam \la0_probe12~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe11~FF  (.D(oTestPort[7]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(la0_probe11)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe11~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe11~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe11~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe11~FF .D_POLARITY = 1'b1;
    defparam \la0_probe11~FF .SR_SYNC = 1'b0;
    defparam \la0_probe11~FF .SR_VALUE = 1'b0;
    defparam \la0_probe11~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe7~FF  (.D(oTestPort[10]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(la0_probe7)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe7~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe7~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe7~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe7~FF .D_POLARITY = 1'b1;
    defparam \la0_probe7~FF .SR_SYNC = 1'b0;
    defparam \la0_probe7~FF .SR_VALUE = 1'b0;
    defparam \la0_probe7~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe14~FF  (.D(oTestPort[24]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(la0_probe14)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe14~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe14~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe14~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe14~FF .D_POLARITY = 1'b1;
    defparam \la0_probe14~FF .SR_SYNC = 1'b0;
    defparam \la0_probe14~FF .SR_VALUE = 1'b0;
    defparam \la0_probe14~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe5[0]~FF  (.D(oTestPort[4]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\la0_probe5[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe5[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe5[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe5[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe5[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe5[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe5[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe5[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe13~FF  (.D(MipiDphyRx1_RX_SKEW_CAL_HS_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(la0_probe13)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe13~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe13~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe13~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe13~FF .D_POLARITY = 1'b1;
    defparam \la0_probe13~FF .SR_SYNC = 1'b0;
    defparam \la0_probe13~FF .SR_VALUE = 1'b0;
    defparam \la0_probe13~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[0]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[0]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\la0_probe6[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe6[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe3~FF  (.D(MipiDphyRx1_ERR_SOT_HS_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(la0_probe3)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe3~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe3~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe3~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe3~FF .D_POLARITY = 1'b1;
    defparam \la0_probe3~FF .SR_SYNC = 1'b0;
    defparam \la0_probe3~FF .SR_VALUE = 1'b0;
    defparam \la0_probe3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9~FF  (.D(MipiDphyRx1_ERR_SOT_SYNC_HS_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(la0_probe9)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe9~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe17~FF  (.D(MipiDphyRx1_STOPSTATE_CLK), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(la0_probe17)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsiRxController.v(361)
    defparam \la0_probe17~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe17~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe17~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe17~FF .D_POLARITY = 1'b1;
    defparam \la0_probe17~FF .SR_SYNC = 1'b0;
    defparam \la0_probe17~FF .SR_VALUE = 1'b0;
    defparam \la0_probe17~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(115)
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wCddFifoFull~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qFullAllmost ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(wCddFifoFull)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(105)
    defparam \wCddFifoFull~FF .CLK_POLARITY = 1'b1;
    defparam \wCddFifoFull~FF .CE_POLARITY = 1'b1;
    defparam \wCddFifoFull~FF .SR_POLARITY = 1'b0;
    defparam \wCddFifoFull~FF .D_POLARITY = 1'b1;
    defparam \wCddFifoFull~FF .SR_SYNC = 1'b0;
    defparam \wCddFifoFull~FF .SR_VALUE = 1'b0;
    defparam \wCddFifoFull~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsValid~FF  (.D(\MCsiRxController/MCsi2Decoder/n640 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsValid )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsValid~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/wHsValid~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsValid~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/select_39/Select_2/n15 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\MCsiRxController/MCsi2Decoder/rHsSt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(226)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/select_39/Select_1/n17 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\MCsiRxController/MCsi2Decoder/rHsSt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(226)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[7]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[6]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[5]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[4]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[3]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[2]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[1]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n21 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/wFtiEmp[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(112)
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_VALUE = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF  (.D(n3753), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF  (.D(n3751), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF  (.D(n3749), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF  (.D(n3747), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF  (.D(n3745), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF  (.D(n3743), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF  (.D(n3741), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF  (.D(n3739), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF  (.D(n3737), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10]_2~FF  (.D(n3736), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n265 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n270 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n275 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n280 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n285 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n290 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n295 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n300 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n305 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n310 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[9] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[10]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[10] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[11]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[11] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[12]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[12] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[13]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[13] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[13]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[14]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[14] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[14]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[15]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[15] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/wHsPixel[15]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[9] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[10] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[11] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[12] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[13] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[14] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[15] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[1] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[10]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[11]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[11]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[12]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[12]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[13]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[13]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[13]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[14]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[6] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[14]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[14]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[15]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[7] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsWordCnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[15]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[15]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsDatatype[2]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[2]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[2]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsDatatype[3]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[3]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[3]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsDatatype[4]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[4]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[4]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \wHsDatatype[5]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[5]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[5]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF  (.D(n129), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF  (.D(n3734), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF  (.D(n3732), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF  (.D(n3730), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF  (.D(n3728), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF  (.D(n3726), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF  (.D(n3724), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF  (.D(n3722), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF  (.D(n3720), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF  (.D(n3718), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF  (.D(n3716), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF  (.D(n3715), 
           .CE(\MCsiRxController/MCsi2Decoder/n659 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(291)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[1]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[2]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[3]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[4]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[5]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[6]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[7]), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wCdcFifoFull_2~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(wCdcFifoFull)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(85)
    defparam \wCdcFifoFull_2~FF .CLK_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .CE_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .SR_POLARITY = 1'b0;
    defparam \wCdcFifoFull_2~FF .D_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .SR_SYNC = 1'b0;
    defparam \wCdcFifoFull_2~FF .SR_VALUE = 1'b0;
    defparam \wCdcFifoFull_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wVideoVd~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/qRVD ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(wVideoVd)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(91)
    defparam \wVideoVd~FF .CLK_POLARITY = 1'b1;
    defparam \wVideoVd~FF .CE_POLARITY = 1'b1;
    defparam \wVideoVd~FF .SR_POLARITY = 1'b0;
    defparam \wVideoVd~FF .D_POLARITY = 1'b1;
    defparam \wVideoVd~FF .SR_SYNC = 1'b0;
    defparam \wVideoVd~FF .SR_VALUE = 1'b0;
    defparam \wVideoVd~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wFtiEmp[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/wFtiEmp[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(88)
    defparam \MCsiRxController/wFtiEmp[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_VALUE = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF  (.D(n106), .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF  (.D(n183), .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF  (.D(n3713), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF  (.D(n3711), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF  (.D(n3709), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF  (.D(n3707), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF  (.D(n3705), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF  (.D(n3704), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n436 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n441 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n446 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n451 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n456 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n461 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n466 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n471 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[0]~FF  (.D(\MVideoPostProcess/rVtgRstCnt[0] ), 
           .CE(\MVideoPostProcess/qVtgRstCntCke ), .CLK(iVCLK), .SR(rVRST), 
           .Q(\MVideoPostProcess/rVtgRstCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[0]~FF  (.D(\MVideoPostProcess/rVtgRstSel ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRST[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstSel_2~FF  (.D(1'b0), .CE(\MVideoPostProcess/equal_18/n21 ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstSel )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n816 ), 
           .CE(\~ceg_net510 ), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n833 ), 
           .CE(\~ceg_net510 ), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_last_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1235 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] ), 
           .CE(ceg_net477), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF  (.D(ceg_net42), 
           .CE(ceg_net1377), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1243 ), .CLK(iBCLK), 
           .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1243 ), .CLK(iBCLK), 
           .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 ), 
           .CE(ceg_net1421), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511SdaOe~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 ), 
           .CE(ceg_net1389), .CLK(iBCLK), .SR(rBRST), .Q(oAdv7511SdaOe)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \oAdv7511SdaOe~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .CE_POLARITY = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .SR_SYNC = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511SclOe~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 ), 
           .CE(ceg_net567), .CLK(iBCLK), .SR(rBRST), .Q(oAdv7511SclOe)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \oAdv7511SclOe~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .CE_POLARITY = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .SR_SYNC = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 ), 
           .CE(ceg_net1523), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 ), 
           .CE(ceg_net1415), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/w_ack~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/w_ack )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 ), 
           .CE(ceg_net617), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0_2~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_0_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 ), 
           .CE(ceg_net1421), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 ), 
           .CE(ceg_net1421), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 ), 
           .CE(ceg_net1460), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 ), 
           .CE(ceg_net1523), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 ), 
           .CE(ceg_net1523), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 ), 
           .CE(ceg_net1523), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 ), 
           .CE(ceg_net1523), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 ), 
           .CE(ceg_net1523), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 ), 
           .CE(ceg_net1523), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 ), 
           .CE(ceg_net1523), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 ), 
           .CE(ceg_net1531), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 ), 
           .CE(ceg_net1415), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 ), 
           .CE(ceg_net1415), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n10449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4687)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n10448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4701)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4  (.I0(n9980), 
            .I1(1'b1), .CI(1'b0), .CO(n10447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4  (.I0(n9781), 
            .I1(1'b1), .CI(1'b0), .CO(n10446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n253 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n252 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n251 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n250 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n249 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n248 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n247 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n246 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n245 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n244 ), 
           .CE(ceg_net941), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n700 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n705 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n710 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n715 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n720 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n725 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n730 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n735 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n740 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n745 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n750 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n755 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n760 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n765 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n770 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n780 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1235 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n785 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1235 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n790 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1235 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n795 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1235 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n800 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1235 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n805 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1235 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n810 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1235 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] ), 
           .CE(ceg_net477), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] ), 
           .CE(ceg_net477), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] ), 
           .CE(ceg_net477), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] ), 
           .CE(ceg_net477), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] ), 
           .CE(ceg_net477), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] ), 
           .CE(ceg_net477), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] ), 
           .CE(ceg_net477), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
           .CE(ceg_net1377), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/sample/adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n131 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rFvde[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/qVde ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rFvde[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511Hs~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rHSync[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511Hs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \oAdv7511Hs~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511Hs~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511Hs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n130 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n129 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF  (.D(n3652), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF  (.D(n3650), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n126 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n125 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF  (.D(n3644), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF  (.D(n3642), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF  (.D(n3640), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n121 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF  (.D(n3637), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511Vs~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVSync[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511Vs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \oAdv7511Vs~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511Vs~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511Vs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511De~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVde[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511De)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(120)
    defparam \oAdv7511De~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511De~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511De~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rFvde[1]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rFvde[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rFvde[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rFvde[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/wVgaGenFDe~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rFvde[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/wVgaGenFDe )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/wVgaGenFDe~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/wVgaGenFDe~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF  (.D(n386), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF  (.D(n3673), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF  (.D(n3671), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF  (.D(n3669), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF  (.D(n3667), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF  (.D(n3665), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF  (.D(n3663), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF  (.D(n3661), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF  (.D(n3659), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF  (.D(n3657), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF  (.D(n3656), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wVideofull~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(wVideofull)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(105)
    defparam \wVideofull~FF .CLK_POLARITY = 1'b1;
    defparam \wVideofull~FF .CE_POLARITY = 1'b1;
    defparam \wVideofull~FF .SR_POLARITY = 1'b0;
    defparam \wVideofull~FF .D_POLARITY = 1'b1;
    defparam \wVideofull~FF .SR_SYNC = 1'b0;
    defparam \wVideofull~FF .SR_VALUE = 1'b0;
    defparam \wVideofull~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n444), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n3635), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3633), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3631), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3629), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3627), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3625), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3623), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3621), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3619), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3617), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3616), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n483 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n488 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n493 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n498 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n503 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n508 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n513 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n518 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n523 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n528 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n533 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n508), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n481), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3614), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3612), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3610), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3608), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3606), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3604), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3602), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3600), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3598), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3597), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n552), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n525), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3595), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3593), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3591), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3589), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3587), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3585), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3583), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3581), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3579), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3578), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n596), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n569), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3576), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3574), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3572), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3570), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3568), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3566), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3564), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3562), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3560), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3559), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n640), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n613), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3557), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3555), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3553), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3551), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3549), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3547), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3545), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3543), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3541), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3540), 
           .CE(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n684), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n657), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3538), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3536), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3534), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3532), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3530), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3528), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3526), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3524), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3522), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3521), 
           .CE(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n728), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n701), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3519), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3517), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3515), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3513), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3511), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3509), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3507), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3505), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3503), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3502), 
           .CE(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n772), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n745), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3500), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3498), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3496), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3494), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3492), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3490), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3488), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3486), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3484), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3483), 
           .CE(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n816), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n789), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3481), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3479), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3477), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3475), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3473), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3471), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3469), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3467), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3465), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3464), 
           .CE(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__13846 (.I0(\MCsiRxController/MCsi2Decoder/wFtiRd[16] ), 
            .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), .I2(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .O(n10054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc1f */ ;
    defparam LUT__13846.LUTMASK = 16'hfc1f;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n860), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n833), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3462), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3460), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3458), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3456), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3454), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3452), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3450), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3448), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3446), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3445), 
           .CE(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n904), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n877), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3443), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3441), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3439), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3437), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3435), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3433), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3431), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3429), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3427), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3426), 
           .CE(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n948), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n921), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3424), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3422), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3420), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3418), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3416), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3414), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3412), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3410), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3408), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3407), 
           .CE(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n992), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n965), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3405), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3403), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3401), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3399), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3397), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3395), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3393), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3391), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3389), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3388), 
           .CE(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n1036), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n1009), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3386), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3384), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3382), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3380), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3378), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3376), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3374), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3372), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3370), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3369), 
           .CE(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n1080), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n1053), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3367), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3365), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3363), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3361), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3359), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3357), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3355), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3353), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3351), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3350), 
           .CE(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RESET_N), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF  (.D(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n1124), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n1097), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n3348), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n3346), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n3344), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n3342), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n3340), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n3338), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n3336), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n3334), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF  (.D(n3332), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF  (.D(n3331), 
           .CE(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[1]~FF  (.D(n268), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[2]~FF  (.D(n304), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[3]~FF  (.D(n3702), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[4]~FF  (.D(n3700), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[5]~FF  (.D(n3698), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[6]~FF  (.D(n3696), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[7]~FF  (.D(n3694), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[8]~FF  (.D(n3692), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[9]~FF  (.D(n3690), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[10]~FF  (.D(n3689), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[1]~FF  (.D(\MVideoPostProcess/rVtgRST[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRST[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[2]_2~FF  (.D(\MVideoPostProcess/rVtgRST[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(183)
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[5]~FF  (.D(oLed[5]), .CE(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), 
           .CLK(iSCLK), .SR(rSRST), .Q(oLed[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(71)
    defparam \oLed[5]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[5]~FF .CE_POLARITY = 1'b0;
    defparam \oLed[5]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[5]~FF .D_POLARITY = 1'b0;
    defparam \oLed[5]~FF .SR_SYNC = 1'b1;
    defparam \oLed[5]~FF .SR_VALUE = 1'b0;
    defparam \oLed[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF  (.D(wVideoVd), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF  (.D(n1167), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF  (.D(n1141), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF  (.D(n3329), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF  (.D(n3327), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF  (.D(n3325), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF  (.D(n3323), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF  (.D(n3321), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF  (.D(n3319), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF  (.D(n3317), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF  (.D(n3315), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF  (.D(n3314), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[1].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[4]~FF  (.D(oLed[4]), .CE(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] ), 
           .CLK(iSCLK), .SR(rSRST), .Q(oLed[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(71)
    defparam \oLed[4]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[4]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[4]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[4]~FF .D_POLARITY = 1'b0;
    defparam \oLed[4]~FF .SR_SYNC = 1'b1;
    defparam \oLed[4]~FF .SR_VALUE = 1'b0;
    defparam \oLed[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF  (.D(wCddFifoFull), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[1].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF  (.D(\genblk1.genblk1[1].mPulseGenerator/n50 ), 
           .CE(\genblk1.genblk1[1].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[1].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[1].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[1].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[1].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[2]~FF  (.D(oLed[2]), .CE(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), 
           .CLK(iSCLK), .SR(rSRST), .Q(oLed[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(71)
    defparam \oLed[2]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[2]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[2]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[2]~FF .D_POLARITY = 1'b0;
    defparam \oLed[2]~FF .SR_SYNC = 1'b1;
    defparam \oLed[2]~FF .SR_VALUE = 1'b0;
    defparam \oLed[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF  (.D(wCdcFifoFull), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/n50 ), 
           .CE(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[1]~FF  (.D(oLed[1]), .CE(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), 
           .CLK(iSCLK), .SR(rSRST), .Q(oLed[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(71)
    defparam \oLed[1]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[1]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[1]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[1]~FF .D_POLARITY = 1'b0;
    defparam \oLed[1]~FF .SR_SYNC = 1'b1;
    defparam \oLed[1]~FF .SR_VALUE = 1'b0;
    defparam \oLed[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF  (.D(wVideofull), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/n50 ), 
           .CE(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 ), .CLK(iSCLK), 
           .SR(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(54)
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n1325 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1326 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1327 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n1950 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3711)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[0] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3740)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n2174 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[0] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2451 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state[0] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3822)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_soft_reset_in ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4132)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2751 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_soft_reset_in ), 
           .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4132)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(la0_probe0), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(la0_probe1), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3584 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF  (.D(la0_probe2), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4417 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF  (.D(la0_probe3), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF  (.D(la0_probe4), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6083 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF  (.D(\la0_probe5[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6972 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6987 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7185 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF  (.D(\la0_probe6[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7869 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7884 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF  (.D(la0_probe7), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8710 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF  (.D(la0_probe8), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9543 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF  (.D(la0_probe9), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10376 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF  (.D(la0_probe10), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n11209 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF  (.D(la0_probe11), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n12042 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF  (.D(la0_probe12), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n12875 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF  (.D(la0_probe13), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n13708 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF  (.D(la0_probe14), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n14541 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF  (.D(la0_probe15), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0]~FF  (.D(la0_probe16), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n16207 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0]~FF  (.D(la0_probe17), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n17040 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0]~FF  (.D(\la0_probe18[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n17887 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n17902 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n18100 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1381 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3684)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1898 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3696)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[1] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[2] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[3] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[4] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[5] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[6] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[7] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[8] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[9] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[10] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[11] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[12] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[13] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[14] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[15] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[16] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[17] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[18] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[19] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[20] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[21] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[22] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[23] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[24] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[25]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[25] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[26]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[26] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[27]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[27] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3730)
    defparam \edb_top_inst/la0/address_counter[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3740)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3740)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3740)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n2173 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n2172 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n2171 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n2170 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n2169 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[1] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[2] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[3] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[4] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[5] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[6] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[7] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[8] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[9] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[10] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[11] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[12] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[13] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[14] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[15] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3767)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2450 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2449 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2448 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2447 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2446 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2445 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2444 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2443 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2442 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2441 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2440 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2439 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2438 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2437 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2436 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2435 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2434 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2433 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2432 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2431 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2430 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2429 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2428 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2427 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2426 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2425 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2424 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2423 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2422 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2421 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2420 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2419 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2418 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2417 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2416 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2415 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2414 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2413 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2412 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2411 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2410 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2409 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2408 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2407 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2406 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2405 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2404 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2403 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2402 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2401 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2400 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2399 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2398 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2397 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2396 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2395 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2394 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2393 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2392 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2391 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2390 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2389 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2388 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3780)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state[1] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3822)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state[2] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3822)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state[3] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3822)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n150 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n149 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n148 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n147 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n146 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n145 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n144 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n143 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n142 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n141 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n140 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n139 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n138 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n137 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n136 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n135 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n134 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n133 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n132 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n131 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n130 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n129 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n128 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n127 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n126 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n125 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n124 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n123 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n122 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n121 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n120 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n119 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(312)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2751 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n2751 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3584 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3584 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4417 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4417 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5250 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6083 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6083 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6972 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6972 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6987 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6987 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n6987 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n6987 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n6987 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n6987 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n6987 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7185 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7185 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n7185 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n7185 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n7185 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n7185 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n7185 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n21 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n20 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7869 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7869 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7884 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7884 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n7884 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n7884 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n7884 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n7884 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n7884 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n8082 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n21 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n20 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8710 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8710 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9543 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9543 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10376 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10376 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n11209 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n11209 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n12042 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n12042 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n12875 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n12875 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n13708 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n13708 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n14541 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n14541 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n15374 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n15374 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n15374 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n16207 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n16207 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n17040 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n17040 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4159)
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5611)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5550)
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n17887 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n17887 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4251)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n17902 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4267)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n18100 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4283)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n10 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/equal_9/n3 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n26 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n9 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5662)
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n131 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5792)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5278)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5078)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5078)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5078)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5314)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5314)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5314)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5324)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5337)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5337)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5337)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5461)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1288 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/n25424 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5278)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5278)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5278)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5078)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n374 ), 
           .CE(\edb_top_inst/ceg_net348 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5349)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF  (.D(\edb_top_inst/la0/address_counter[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF  (.D(\edb_top_inst/la0/address_counter[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[27]~FF  (.D(\edb_top_inst/la0/address_counter[27] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n374 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5359)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[1] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[2] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[5] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[6] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[7] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[8] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[9] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[10] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[11] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[12] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[13]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[13] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[14]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[14] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[15]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[16]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[17]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[18]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[19]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[20]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[21]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[22]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[23]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[24]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[25]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[26]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[27]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[27] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[28]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[28] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[29]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[29] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[30]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[30] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[31]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[31] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[32]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[32] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[33]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[33] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[34]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[34] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1303 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5368)
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5461)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/n2043 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/n1019 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/n1017 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/n1015 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/n1013 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/n1011 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/n1009 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/n1007 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/n1005 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/n1003 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF  (.D(\edb_top_inst/n1001 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF  (.D(\edb_top_inst/n999 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12]~FF  (.D(\edb_top_inst/n998 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/n662 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/n996 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/n994 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/n992 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/n990 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/n988 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/n986 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/n984 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/n981 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF  (.D(\edb_top_inst/n978 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF  (.D(\edb_top_inst/n976 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12]~FF  (.D(\edb_top_inst/n974 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2043 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/n664 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/n971 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/n969 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/n967 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/n965 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/n963 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/n961 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/n959 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/n957 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF  (.D(\edb_top_inst/n955 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF  (.D(\edb_top_inst/n953 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12]~FF  (.D(\edb_top_inst/n951 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/n877 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/n900 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/n898 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/n896 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/n894 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/n892 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/n890 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/n888 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/n886 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/n884 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[11]~FF  (.D(\edb_top_inst/n882 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[12]~FF  (.D(\edb_top_inst/n880 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[13]~FF  (.D(\edb_top_inst/n879 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4708)
    defparam \edb_top_inst/la0/la_sample_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4777)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[12] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[12] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4599)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/n878 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/n923 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/n921 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/n919 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/n917 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/n915 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/n913 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/n911 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/n909 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF  (.D(\edb_top_inst/n907 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF  (.D(\edb_top_inst/n905 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[12]~FF  (.D(\edb_top_inst/n903 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13]~FF  (.D(\edb_top_inst/n902 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4694)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3625)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1297 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3674)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(383)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]_2~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(383)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(383)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(383)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]_2~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]_2~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]_2~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]_2~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]_2~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]_2~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]_2~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]_2~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]_2~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]_2~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]_2~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]_2~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]_2~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]_2~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]_2~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]_2~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]_2~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]_2~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]_2~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]_2~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]_2~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]_2~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]_2~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]_2~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]_2~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]_2~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]_2~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]_2~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]_2~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]_2~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]_2~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]_2~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]_2~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]_2~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]_2~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]_2~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]_2~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]_2~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]_2~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]_2~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]_2~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]_2~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]_2~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]_2~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]_2~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]_2~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]_2~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]_2~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]_2~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]_2~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]_2~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]_2~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]_2~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]_2~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]_2~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]_2~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]_2~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]_2~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]_2~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]_2~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]_2~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]_2~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]_2~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]_2~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]_2~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]_2~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]_2~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]_2~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]_2~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]_2~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]_2~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]_2~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]_2~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]_2~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]_2~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]_2~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]_2~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]_2~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]_2~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]_2~FF  (.D(\edb_top_inst/edb_user_dr[81] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]_2~FF  (.D(jtag_inst2_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(376)
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), .CI(1'b0), 
            .O(n106), .CO(n107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i2  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), .CI(1'b0), 
            .O(n129), .CO(n130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n107), .O(n183), .CO(n184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i2  (.I0(\MVideoPostProcess/rVtgRstCnt[1] ), 
            .I1(\MVideoPostProcess/rVtgRstCnt[0] ), .CI(1'b0), .O(n268), 
            .CO(n269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i3  (.I0(\MVideoPostProcess/rVtgRstCnt[2] ), 
            .I1(1'b0), .CI(n269), .O(n304), .CO(n305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i2  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[1] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), .CI(1'b0), 
            .O(n386), .CO(n387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i2  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[1] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), .CI(1'b0), 
            .O(n441), .CO(n442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n444), .CO(n445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n509), .O(n481), .CO(n482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n508), .CO(n509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n553), .O(n525), .CO(n526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n552), .CO(n553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n597), .O(n569), .CO(n570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n596), .CO(n597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n641), .O(n613), .CO(n614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n640), .CO(n641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n685), .O(n657), .CO(n658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n684), .CO(n685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n729), .O(n701), .CO(n702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n728), .CO(n729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n773), .O(n745), .CO(n746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n772), .CO(n773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n817), .O(n789), .CO(n790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n816), .CO(n817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n861), .O(n833), .CO(n834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n860), .CO(n861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n905), .O(n877), .CO(n878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n904), .CO(n905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n949), .O(n921), .CO(n922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n948), .CO(n949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n993), .O(n965), .CO(n966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n992), .CO(n993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n1037), .O(n1009), .CO(n1010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n1036), .CO(n1037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n1081), .O(n1053), .CO(n1054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n1080), .CO(n1081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n1125), .O(n1097), .CO(n1098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n1124), .CO(n1125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i3  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[2] ), 
            .I1(1'b0), .CI(n1168), .O(n1141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i3 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i2  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), .CI(1'b0), 
            .O(n1167), .CO(n1168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i2 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i12  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] ), 
            .I1(1'b0), .CI(n3316), .O(n3314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i12 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i11  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] ), 
            .I1(1'b0), .CI(n3318), .O(n3315), .CO(n3316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i11 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i10  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] ), 
            .I1(1'b0), .CI(n3320), .O(n3317), .CO(n3318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i10 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i9  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] ), 
            .I1(1'b0), .CI(n3322), .O(n3319), .CO(n3320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i9 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i8  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] ), 
            .I1(1'b0), .CI(n3324), .O(n3321), .CO(n3322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i8 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i7  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] ), 
            .I1(1'b0), .CI(n3326), .O(n3323), .CO(n3324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i7 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i6  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] ), 
            .I1(1'b0), .CI(n3328), .O(n3325), .CO(n3326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i6 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i5  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] ), 
            .I1(1'b0), .CI(n3330), .O(n3327), .CO(n3328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i5 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i4  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] ), 
            .I1(1'b0), .CI(n10446), .O(n3329), .CO(n3330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3333), .O(n3331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3335), .O(n3332), .CO(n3333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3337), .O(n3334), .CO(n3335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3339), .O(n3336), .CO(n3337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3341), .O(n3338), .CO(n3339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3343), .O(n3340), .CO(n3341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3345), .O(n3342), .CO(n3343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3347), .O(n3344), .CO(n3345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3349), .O(n3346), .CO(n3347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n1098), .O(n3348), .CO(n3349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3352), .O(n3350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3354), .O(n3351), .CO(n3352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3356), .O(n3353), .CO(n3354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3358), .O(n3355), .CO(n3356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3360), .O(n3357), .CO(n3358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3362), .O(n3359), .CO(n3360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3364), .O(n3361), .CO(n3362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3366), .O(n3363), .CO(n3364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3368), .O(n3365), .CO(n3366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n1054), .O(n3367), .CO(n3368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3371), .O(n3369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3373), .O(n3370), .CO(n3371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3375), .O(n3372), .CO(n3373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3377), .O(n3374), .CO(n3375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3379), .O(n3376), .CO(n3377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3381), .O(n3378), .CO(n3379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3383), .O(n3380), .CO(n3381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3385), .O(n3382), .CO(n3383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3387), .O(n3384), .CO(n3385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n1010), .O(n3386), .CO(n3387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3390), .O(n3388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3392), .O(n3389), .CO(n3390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3394), .O(n3391), .CO(n3392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3396), .O(n3393), .CO(n3394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3398), .O(n3395), .CO(n3396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3400), .O(n3397), .CO(n3398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3402), .O(n3399), .CO(n3400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3404), .O(n3401), .CO(n3402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3406), .O(n3403), .CO(n3404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n966), .O(n3405), .CO(n3406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3409), .O(n3407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3411), .O(n3408), .CO(n3409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3413), .O(n3410), .CO(n3411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3415), .O(n3412), .CO(n3413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3417), .O(n3414), .CO(n3415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3419), .O(n3416), .CO(n3417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3421), .O(n3418), .CO(n3419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3423), .O(n3420), .CO(n3421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3425), .O(n3422), .CO(n3423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n922), .O(n3424), .CO(n3425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3428), .O(n3426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3430), .O(n3427), .CO(n3428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3432), .O(n3429), .CO(n3430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3434), .O(n3431), .CO(n3432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3436), .O(n3433), .CO(n3434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3438), .O(n3435), .CO(n3436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3440), .O(n3437), .CO(n3438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3442), .O(n3439), .CO(n3440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3444), .O(n3441), .CO(n3442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n878), .O(n3443), .CO(n3444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3447), .O(n3445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3449), .O(n3446), .CO(n3447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3451), .O(n3448), .CO(n3449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3453), .O(n3450), .CO(n3451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3455), .O(n3452), .CO(n3453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3457), .O(n3454), .CO(n3455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3459), .O(n3456), .CO(n3457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3461), .O(n3458), .CO(n3459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3463), .O(n3460), .CO(n3461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n834), .O(n3462), .CO(n3463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3466), .O(n3464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3468), .O(n3465), .CO(n3466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3470), .O(n3467), .CO(n3468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3472), .O(n3469), .CO(n3470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3474), .O(n3471), .CO(n3472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3476), .O(n3473), .CO(n3474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3478), .O(n3475), .CO(n3476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3480), .O(n3477), .CO(n3478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3482), .O(n3479), .CO(n3480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n790), .O(n3481), .CO(n3482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3485), .O(n3483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3487), .O(n3484), .CO(n3485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3489), .O(n3486), .CO(n3487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3491), .O(n3488), .CO(n3489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3493), .O(n3490), .CO(n3491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3495), .O(n3492), .CO(n3493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3497), .O(n3494), .CO(n3495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3499), .O(n3496), .CO(n3497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3501), .O(n3498), .CO(n3499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n746), .O(n3500), .CO(n3501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3504), .O(n3502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3506), .O(n3503), .CO(n3504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3508), .O(n3505), .CO(n3506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3510), .O(n3507), .CO(n3508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3512), .O(n3509), .CO(n3510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3514), .O(n3511), .CO(n3512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3516), .O(n3513), .CO(n3514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3518), .O(n3515), .CO(n3516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3520), .O(n3517), .CO(n3518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n702), .O(n3519), .CO(n3520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3523), .O(n3521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3525), .O(n3522), .CO(n3523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3527), .O(n3524), .CO(n3525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3529), .O(n3526), .CO(n3527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3531), .O(n3528), .CO(n3529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3533), .O(n3530), .CO(n3531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3535), .O(n3532), .CO(n3533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3537), .O(n3534), .CO(n3535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3539), .O(n3536), .CO(n3537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n658), .O(n3538), .CO(n3539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3542), .O(n3540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3544), .O(n3541), .CO(n3542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3546), .O(n3543), .CO(n3544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3548), .O(n3545), .CO(n3546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3550), .O(n3547), .CO(n3548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3552), .O(n3549), .CO(n3550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3554), .O(n3551), .CO(n3552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3556), .O(n3553), .CO(n3554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3558), .O(n3555), .CO(n3556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n614), .O(n3557), .CO(n3558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3561), .O(n3559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3563), .O(n3560), .CO(n3561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3565), .O(n3562), .CO(n3563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3567), .O(n3564), .CO(n3565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3569), .O(n3566), .CO(n3567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3571), .O(n3568), .CO(n3569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3573), .O(n3570), .CO(n3571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3575), .O(n3572), .CO(n3573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3577), .O(n3574), .CO(n3575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n570), .O(n3576), .CO(n3577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3580), .O(n3578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3582), .O(n3579), .CO(n3580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3584), .O(n3581), .CO(n3582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3586), .O(n3583), .CO(n3584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3588), .O(n3585), .CO(n3586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3590), .O(n3587), .CO(n3588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3592), .O(n3589), .CO(n3590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3594), .O(n3591), .CO(n3592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3596), .O(n3593), .CO(n3594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n526), .O(n3595), .CO(n3596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3599), .O(n3597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3601), .O(n3598), .CO(n3599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3603), .O(n3600), .CO(n3601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3605), .O(n3602), .CO(n3603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3607), .O(n3604), .CO(n3605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3609), .O(n3606), .CO(n3607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3611), .O(n3608), .CO(n3609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3613), .O(n3610), .CO(n3611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3615), .O(n3612), .CO(n3613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n482), .O(n3614), .CO(n3615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i13  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
            .I1(1'b0), .CI(n3618), .O(n3616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i13 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i12  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
            .I1(1'b0), .CI(n3620), .O(n3617), .CO(n3618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n3622), .O(n3619), .CO(n3620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n3624), .O(n3621), .CO(n3622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3626), .O(n3623), .CO(n3624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3628), .O(n3625), .CO(n3626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3630), .O(n3627), .CO(n3628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3632), .O(n3629), .CO(n3630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3634), .O(n3631), .CO(n3632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n3636), .O(n3633), .CO(n3634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n445), .O(n3635), .CO(n3636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i12  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I1(1'b0), .CI(n3639), .O(n3637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i11  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I1(1'b0), .CI(n3641), .O(n3638), .CO(n3639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i10  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[9] ), 
            .I1(1'b0), .CI(n3643), .O(n3640), .CO(n3641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i9  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[8] ), 
            .I1(1'b0), .CI(n3645), .O(n3642), .CO(n3643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i8  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[7] ), 
            .I1(1'b0), .CI(n3647), .O(n3644), .CO(n3645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i7  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), 
            .I1(1'b0), .CI(n3649), .O(n3646), .CO(n3647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i6  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), 
            .I1(1'b0), .CI(n3651), .O(n3648), .CO(n3649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i5  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I1(1'b0), .CI(n3653), .O(n3650), .CO(n3651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i4  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .I1(1'b0), .CI(n3655), .O(n3652), .CO(n3653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i3  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .I1(1'b0), .CI(n442), .O(n3654), .CO(n3655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i12  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), 
            .I1(1'b0), .CI(n3658), .O(n3656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i11  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), 
            .I1(1'b0), .CI(n3660), .O(n3657), .CO(n3658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i10  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), 
            .I1(1'b0), .CI(n3662), .O(n3659), .CO(n3660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i9  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), 
            .I1(1'b0), .CI(n3664), .O(n3661), .CO(n3662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i8  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I1(1'b0), .CI(n3666), .O(n3663), .CO(n3664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i7  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I1(1'b0), .CI(n3668), .O(n3665), .CO(n3666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i6  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), 
            .I1(1'b0), .CI(n3670), .O(n3667), .CO(n3668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i5  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), 
            .I1(1'b0), .CI(n3672), .O(n3669), .CO(n3670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i4  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), 
            .I1(1'b0), .CI(n10447), .O(n3671), .CO(n3672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i3  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .I1(1'b0), .CI(n387), .O(n3673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i11  (.I0(\MVideoPostProcess/rVtgRstCnt[10] ), 
            .I1(1'b0), .CI(n3691), .O(n3689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i10  (.I0(\MVideoPostProcess/rVtgRstCnt[9] ), 
            .I1(1'b0), .CI(n3693), .O(n3690), .CO(n3691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i9  (.I0(\MVideoPostProcess/rVtgRstCnt[8] ), 
            .I1(1'b0), .CI(n3695), .O(n3692), .CO(n3693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i8  (.I0(\MVideoPostProcess/rVtgRstCnt[7] ), 
            .I1(1'b0), .CI(n3697), .O(n3694), .CO(n3695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i7  (.I0(\MVideoPostProcess/rVtgRstCnt[6] ), 
            .I1(1'b0), .CI(n3699), .O(n3696), .CO(n3697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i6  (.I0(\MVideoPostProcess/rVtgRstCnt[5] ), 
            .I1(1'b0), .CI(n3701), .O(n3698), .CO(n3699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i5  (.I0(\MVideoPostProcess/rVtgRstCnt[4] ), 
            .I1(1'b0), .CI(n3703), .O(n3700), .CO(n3701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i4  (.I0(\MVideoPostProcess/rVtgRstCnt[3] ), 
            .I1(1'b0), .CI(n305), .O(n3702), .CO(n3703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MVideoPostProcess/MVideoPostProcess.v(169)
    defparam \MVideoPostProcess/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n3706), .O(n3704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n3708), .O(n3705), .CO(n3706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n3710), .O(n3707), .CO(n3708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n3712), .O(n3709), .CO(n3710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n3714), .O(n3711), .CO(n3712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n184), .O(n3713), .CO(n3714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i13  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] ), 
            .I1(1'b0), .CI(n3717), .O(n3715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i13 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i12  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .I1(1'b0), .CI(n3719), .O(n3716), .CO(n3717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i12 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i11  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I1(1'b0), .CI(n3721), .O(n3718), .CO(n3719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i11 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i10  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] ), 
            .I1(1'b0), .CI(n3723), .O(n3720), .CO(n3721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i9  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] ), 
            .I1(1'b0), .CI(n3725), .O(n3722), .CO(n3723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i8  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] ), 
            .I1(1'b0), .CI(n3727), .O(n3724), .CO(n3725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i7  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] ), 
            .I1(1'b0), .CI(n3729), .O(n3726), .CO(n3727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i6  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] ), 
            .I1(1'b0), .CI(n3731), .O(n3728), .CO(n3729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i5  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] ), 
            .I1(1'b0), .CI(n3733), .O(n3730), .CO(n3731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i4  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] ), 
            .I1(1'b0), .CI(n3735), .O(n3732), .CO(n3733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_64/i3  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] ), 
            .I1(1'b0), .CI(n130), .O(n3734), .CO(n3735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/MCsiRxController/MCsi2Decoder.v(287)
    defparam \MCsiRxController/MCsi2Decoder/add_64/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_64/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i11  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10] ), 
            .I1(1'b0), .CI(n3738), .O(n3736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I1(1'b0), .CI(n3740), .O(n3737), .CO(n3738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(1'b0), .CI(n3742), .O(n3739), .CO(n3740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(1'b0), .CI(n3744), .O(n3741), .CO(n3742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(1'b0), .CI(n3746), .O(n3743), .CO(n3744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I1(1'b0), .CI(n3748), .O(n3745), .CO(n3746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(1'b0), .CI(n3750), .O(n3747), .CO(n3748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(1'b0), .CI(n3752), .O(n3749), .CO(n3750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(1'b0), .CI(n3754), .O(n3751), .CO(n3752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .CI(1'b0), .O(n3753), .CO(n3754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/src/common/fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_RAM10 \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2  (.WCLK(oTestPort[17]), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd }), 
            .WDATA({\MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[4] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[3] , 
            \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[2] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[1] , 
            \la0_probe6[0] }), .WADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] }), 
            .RADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] }), 
            .RDATA({\MCsiRxController/MCsi2Decoder/wFtiRd[4] , \MCsiRxController/MCsi2Decoder/wFtiRd[3] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[2] , \MCsiRxController/MCsi2Decoder/wFtiRd[1] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .READ_WIDTH = 5;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .WRITE_WIDTH = 5;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .RESET_OUTREG = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .OUTPUT_REG = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .WRITE_MODE = "READ_UNKNOWN";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$2 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12  (.WCLK(oTestPort[17]), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd }), 
            .WDATA({\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[1] , \la0_probe5[0] , 
            \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[7] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[6] , 
            \MCsiRxController/MCsi2Decoder/rDphyHsDataLane0[5] }), .WADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] }), 
            .RADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] }), 
            .RDATA({\MCsiRxController/MCsi2Decoder/wFtiRd[9] , \MCsiRxController/MCsi2Decoder/wFtiRd[8] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[7] , \MCsiRxController/MCsi2Decoder/wFtiRd[6] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .READ_WIDTH = 5;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .WRITE_WIDTH = 5;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .RESET_OUTREG = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .OUTPUT_REG = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .WRITE_MODE = "READ_UNKNOWN";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12  (.WCLK(oTestPort[17]), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd }), 
            .WDATA({\MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[6] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[5] , 
            \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[4] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[3] , 
            \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[2] }), .WADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] }), 
            .RADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] }), 
            .RDATA({\MCsiRxController/MCsi2Decoder/wFtiRd[14] , \MCsiRxController/MCsi2Decoder/wFtiRd[13] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[12] , \MCsiRxController/MCsi2Decoder/wFtiRd[11] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .READ_WIDTH = 5;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .WRITE_WIDTH = 5;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .RESET_OUTREG = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .OUTPUT_REG = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .WRITE_MODE = "READ_UNKNOWN";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$b12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1  (.WCLK(oTestPort[17]), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd }), 
            .WDATA({3'b000, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs , 
            \MCsiRxController/MCsi2Decoder/rDphyHsDataLane1[7] }), .WADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] }), 
            .RADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] }), 
            .RDATA({Open_0, Open_1, Open_2, \MCsiRxController/MCsi2Decoder/wFtiRd[16] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[15] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=5, WRITE_WIDTH=5, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .READ_WIDTH = 5;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .WRITE_WIDTH = 5;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .RESET_OUTREG = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .OUTPUT_REG = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .WRITE_MODE = "READ_UNKNOWN";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo__D$c1 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo  (.WCLK(iSCLK), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({\MCsiRxController/wHsValid , \MCsiRxController/wHsValid }), 
            .WDATA({\MCsiRxController/wHsPixel[15] , \MCsiRxController/wHsPixel[14] , 
            \MCsiRxController/wHsPixel[13] , \MCsiRxController/wHsPixel[12] , 
            \MCsiRxController/wHsPixel[11] , \MCsiRxController/wHsPixel[10] , 
            \MCsiRxController/wHsPixel[9] , \MCsiRxController/wHsPixel[8] , 
            \MCsiRxController/wHsPixel[7] , \MCsiRxController/wHsPixel[6] , 
            \MCsiRxController/wHsPixel[5] , \MCsiRxController/wHsPixel[4] , 
            \MCsiRxController/wHsPixel[3] , \MCsiRxController/wHsPixel[2] , 
            \MCsiRxController/wHsPixel[1] , \MCsiRxController/wHsPixel[0] }), 
            .WADDR({\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] }), .RADDR({\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] }), 
            .RDATA({\wVideoPixel[15] , \wVideoPixel[14] , \wVideoPixel[13] , 
            \wVideoPixel[12] , \wVideoPixel[11] , \wVideoPixel[10] , \wVideoPixel[9] , 
            \wVideoPixel[8] , \wVideoPixel[7] , \wVideoPixel[6] , \wVideoPixel[5] , 
            \wVideoPixel[4] , \wVideoPixel[3] , \wVideoPixel[2] , \wVideoPixel[1] , 
            \wVideoPixel[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="NONE", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .READ_WIDTH = 16;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WRITE_WIDTH = 16;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RESET_OUTREG = "NONE";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .OUTPUT_REG = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WRITE_MODE = "READ_FIRST";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_SRL8 \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2  (.D(\MVideoPostProcess/mVideoTimingGen/qVrange ), 
            .CLK(iVCLK), .CE(1'b1), .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1 */ ;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .INIT = 8'h0;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \MVideoPostProcess/mVideoTimingGen/dff_41/i4_2  (.D(\MVideoPostProcess/mVideoTimingGen/qVde ), 
            .CLK(iVCLK), .CE(1'b1), .Q(\MVideoPostProcess/mVideoTimingGen/dff_41/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1 */ ;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_41/i4_2 .INIT = 8'h0;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_41/i4_2 .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_41/i4_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2  (.D(\MVideoPostProcess/mVideoTimingGen/qHrange ), 
            .CLK(iVCLK), .CE(1'b1), .Q(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1 */ ;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .INIT = 8'h0;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .CE_POLARITY = 1'b1;
    EFX_RAM10 \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[0] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[8]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[1] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[9]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[2] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[10]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[3] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[11]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[4] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[12]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[5] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[13]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[6] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[14]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[7] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[15]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[8] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[0]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[9] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[1]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[10] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[2]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[11] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[3]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[12] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[4]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[13] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[5]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[14] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[6]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[15] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[12] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[11] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[7]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_LUT4 \edb_top_inst/LUT__4317  (.I0(\edb_top_inst/la0/crc_data_out[21] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n3116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4317 .LUTMASK = 16'h9009;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[32] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$F12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[33] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$G12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2  (.D(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2  (.D(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i6_2  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i6_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i6_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i6_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i6_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i7_2  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i7_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i7_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i7_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i7_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i1_2  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i1_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i1_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i1_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i1_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i2_2  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i2_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i2_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i2_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i2_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i24_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i24_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i24_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i24_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i24_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2  (.D(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2  (.D(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2  (.D(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i3_2  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i3_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i3_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i3_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i3_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2  (.D(\edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2  (.D(\edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2  (.D(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .CE_POLARITY = 1'b1;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[34] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$H1 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[31] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$E12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[30] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$D12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[29] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$C12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[28] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$B12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[27] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$A12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[26] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$z12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[25] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$y12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[24] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$x12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[23] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$w12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[22] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$v12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[21] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[20] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[19] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[18] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[8] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[9] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[11] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[12] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[13] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[14] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[15] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[16] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[17] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_LUT4 \edb_top_inst/LUT__4318  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/edb_user_dr[67] ), .I2(\edb_top_inst/la0/crc_data_out[18] ), 
            .I3(\edb_top_inst/edb_user_dr[68] ), .O(\edb_top_inst/n3117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4318 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4319  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/edb_user_dr[69] ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .I3(\edb_top_inst/edb_user_dr[70] ), .O(\edb_top_inst/n3118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4319 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4320  (.I0(\edb_top_inst/n3115 ), .I1(\edb_top_inst/n3116 ), 
            .I2(\edb_top_inst/n3117 ), .I3(\edb_top_inst/n3118 ), .O(\edb_top_inst/n3119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4320 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4321  (.I0(\edb_top_inst/la0/crc_data_out[27] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .I3(\edb_top_inst/edb_user_dr[78] ), .O(\edb_top_inst/n3120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4321 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4322  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/edb_user_dr[79] ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n3121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4322 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4323  (.I0(\edb_top_inst/la0/crc_data_out[24] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .I3(\edb_top_inst/edb_user_dr[81] ), .O(\edb_top_inst/n3122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4323 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4324  (.I0(\edb_top_inst/la0/crc_data_out[25] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/la0/crc_data_out[26] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n3123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4324 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4325  (.I0(\edb_top_inst/n3120 ), .I1(\edb_top_inst/n3121 ), 
            .I2(\edb_top_inst/n3122 ), .I3(\edb_top_inst/n3123 ), .O(\edb_top_inst/n3124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4325 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4326  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/edb_user_dr[62] ), .I2(\edb_top_inst/la0/crc_data_out[13] ), 
            .I3(\edb_top_inst/edb_user_dr[63] ), .O(\edb_top_inst/n3125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4326 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4327  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/edb_user_dr[57] ), .I2(\edb_top_inst/la0/crc_data_out[14] ), 
            .I3(\edb_top_inst/edb_user_dr[64] ), .O(\edb_top_inst/n3126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4327 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4328  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/edb_user_dr[58] ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .I3(\edb_top_inst/edb_user_dr[59] ), .O(\edb_top_inst/n3127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4328 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4329  (.I0(\edb_top_inst/la0/crc_data_out[10] ), 
            .I1(\edb_top_inst/edb_user_dr[60] ), .I2(\edb_top_inst/la0/crc_data_out[11] ), 
            .I3(\edb_top_inst/edb_user_dr[61] ), .O(\edb_top_inst/n3128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4329 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4330  (.I0(\edb_top_inst/n3125 ), .I1(\edb_top_inst/n3126 ), 
            .I2(\edb_top_inst/n3127 ), .I3(\edb_top_inst/n3128 ), .O(\edb_top_inst/n3129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4330 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4331  (.I0(\edb_top_inst/la0/crc_data_out[0] ), 
            .I1(\edb_top_inst/edb_user_dr[50] ), .I2(\edb_top_inst/la0/crc_data_out[1] ), 
            .I3(\edb_top_inst/edb_user_dr[51] ), .O(\edb_top_inst/n3130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4331 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4332  (.I0(\edb_top_inst/la0/crc_data_out[6] ), 
            .I1(\edb_top_inst/edb_user_dr[56] ), .I2(\edb_top_inst/la0/crc_data_out[15] ), 
            .I3(\edb_top_inst/edb_user_dr[65] ), .O(\edb_top_inst/n3131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4332 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4333  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/edb_user_dr[54] ), .I2(\edb_top_inst/la0/crc_data_out[5] ), 
            .I3(\edb_top_inst/edb_user_dr[55] ), .O(\edb_top_inst/n3132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4333 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4334  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/edb_user_dr[52] ), .I2(\edb_top_inst/la0/crc_data_out[3] ), 
            .I3(\edb_top_inst/edb_user_dr[53] ), .O(\edb_top_inst/n3133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4334 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4335  (.I0(\edb_top_inst/n3130 ), .I1(\edb_top_inst/n3131 ), 
            .I2(\edb_top_inst/n3132 ), .I3(\edb_top_inst/n3133 ), .O(\edb_top_inst/n3134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4335 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4336  (.I0(\edb_top_inst/n3119 ), .I1(\edb_top_inst/n3124 ), 
            .I2(\edb_top_inst/n3129 ), .I3(\edb_top_inst/n3134 ), .O(\edb_top_inst/n3135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4336 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4337  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n3136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4337 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4338  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[6] ), 
            .I3(\edb_top_inst/la0/word_count[7] ), .O(\edb_top_inst/n3137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4338 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4339  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/la0/word_count[11] ), .I2(\edb_top_inst/la0/word_count[12] ), 
            .I3(\edb_top_inst/la0/word_count[13] ), .O(\edb_top_inst/n3138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4339 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4340  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/la0/word_count[9] ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/la0/word_count[15] ), .O(\edb_top_inst/n3139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4340 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4341  (.I0(\edb_top_inst/n3136 ), .I1(\edb_top_inst/n3137 ), 
            .I2(\edb_top_inst/n3138 ), .I3(\edb_top_inst/n3139 ), .O(\edb_top_inst/n3140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4341 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4342  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/la0/bit_count[2] ), 
            .O(\edb_top_inst/n3141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4342 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4343  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(\edb_top_inst/la0/bit_count[4] ), .I2(\edb_top_inst/la0/bit_count[5] ), 
            .I3(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n3142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4343 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4344  (.I0(\edb_top_inst/n3142 ), .I1(\edb_top_inst/n3141 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n3143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4344 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4345  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n3144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4345 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4346  (.I0(\edb_top_inst/n3140 ), .I1(\edb_top_inst/la0/module_state[1] ), 
            .I2(\edb_top_inst/n3143 ), .I3(\edb_top_inst/n3144 ), .O(\edb_top_inst/n3145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4346 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__4347  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n3146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4347 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4348  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n3147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4348 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__4349  (.I0(\edb_top_inst/n3146 ), .I1(\edb_top_inst/n3145 ), 
            .I2(\edb_top_inst/n3147 ), .O(\edb_top_inst/n3148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4349 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4350  (.I0(\edb_top_inst/n3135 ), .I1(\edb_top_inst/la0/crc_data_out[0] ), 
            .I2(\edb_top_inst/n3148 ), .O(\edb_top_inst/n3149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4350 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4351  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), .I2(\edb_top_inst/n3148 ), 
            .O(\edb_top_inst/n3150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4351 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4352  (.I0(\edb_top_inst/la0/opcode[3] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n3093 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4352 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4353  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n3090 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4353 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4354  (.I0(\edb_top_inst/n3093 ), .I1(\edb_top_inst/la0/bit_count[5] ), 
            .I2(\edb_top_inst/n3090 ), .I3(\edb_top_inst/la0/bit_count[4] ), 
            .O(\edb_top_inst/n3151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4354 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__4355  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n3152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4355 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__4356  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/la0/bit_count[2] ), 
            .I3(\edb_top_inst/n3152 ), .O(\edb_top_inst/n3153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4356 .LUTMASK = 16'hfe7f;
    EFX_LUT4 \edb_top_inst/LUT__4357  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n3154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4357 .LUTMASK = 16'hfe3f;
    EFX_LUT4 \edb_top_inst/LUT__4358  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(\edb_top_inst/n3154 ), .O(\edb_top_inst/n3155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4358 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4359  (.I0(\edb_top_inst/n3151 ), .I1(\edb_top_inst/n3153 ), 
            .I2(\edb_top_inst/n3155 ), .I3(\edb_top_inst/n3140 ), .O(\edb_top_inst/n3156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4359 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4360  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg[1] ), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg[2] ), .I2(\edb_top_inst/debug_hub_inst/module_id_reg[3] ), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg[0] ), .O(\edb_top_inst/n3157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4360 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4361  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n3158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4361 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4362  (.I0(\edb_top_inst/n3158 ), .I1(\edb_top_inst/edb_user_dr[81] ), 
            .I2(\edb_top_inst/n3157 ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n3159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4362 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__4363  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/n3156 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n3159 ), 
            .O(\edb_top_inst/n3160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4363 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__4364  (.I0(jtag_inst2_CAPTURE), .I1(\edb_top_inst/n3157 ), 
            .O(\edb_top_inst/n3161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4364 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4365  (.I0(\edb_top_inst/n3161 ), .I1(\edb_top_inst/n3140 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n3162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4365 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4366  (.I0(\edb_top_inst/n3158 ), .I1(\edb_top_inst/n3156 ), 
            .I2(\edb_top_inst/n3162 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n3163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4366 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4367  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/biu_ready ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n3164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4367 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__4368  (.I0(\edb_top_inst/n3161 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/n3164 ), 
            .O(\edb_top_inst/n3165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4368 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__4369  (.I0(\edb_top_inst/edb_user_dr[77] ), 
            .I1(\edb_top_inst/edb_user_dr[78] ), .I2(\edb_top_inst/edb_user_dr[79] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n3166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4369 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__4370  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(jtag_inst2_UPDATE), .I2(\edb_top_inst/n3157 ), .O(\edb_top_inst/n3167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4370 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4371  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n3168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4371 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4372  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3167 ), 
            .I2(\edb_top_inst/n3168 ), .O(\edb_top_inst/n3169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4372 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4373  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n3165 ), .I2(\edb_top_inst/n3169 ), .O(\edb_top_inst/n3170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4373 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4374  (.I0(\edb_top_inst/n3145 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n3171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4374 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4375  (.I0(\edb_top_inst/n3160 ), .I1(\edb_top_inst/n3163 ), 
            .I2(\edb_top_inst/n3170 ), .I3(\edb_top_inst/n3171 ), .O(\edb_top_inst/la0/module_next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4375 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4376  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n3172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4376 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4377  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4377 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4378  (.I0(\edb_top_inst/la0/module_next_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/n3172 ), 
            .I3(\edb_top_inst/n3173 ), .O(\edb_top_inst/n3174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4378 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__4379  (.I0(\edb_top_inst/n3150 ), .I1(\edb_top_inst/n3149 ), 
            .I2(\edb_top_inst/n3174 ), .I3(\edb_top_inst/n3157 ), .O(jtag_inst2_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4379 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4380  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[40] ), .O(\edb_top_inst/la0/n1325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4380 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4381  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/edb_user_dr[75] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n3175 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4381 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4382  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/edb_user_dr[68] ), .I2(\edb_top_inst/edb_user_dr[69] ), 
            .I3(\edb_top_inst/edb_user_dr[79] ), .O(\edb_top_inst/n3176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4382 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4383  (.I0(\edb_top_inst/edb_user_dr[78] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/edb_user_dr[80] ), 
            .O(\edb_top_inst/n3177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4383 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4384  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n3168 ), .O(\edb_top_inst/n3178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4384 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4385  (.I0(\edb_top_inst/n3167 ), .I1(\edb_top_inst/n3176 ), 
            .I2(\edb_top_inst/n3177 ), .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/n3179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4385 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4386  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n3179 ), .O(\edb_top_inst/n3180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4386 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4387  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n3180 ), 
            .O(\edb_top_inst/n3181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4387 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4388  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .I3(\edb_top_inst/n3181 ), .O(\edb_top_inst/n3182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4388 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4389  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/n3175 ), 
            .I2(\edb_top_inst/la0/la_soft_reset_in ), .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4389 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4390  (.I0(\edb_top_inst/n3175 ), .I1(\edb_top_inst/n3182 ), 
            .O(\edb_top_inst/la0/n1297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4390 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4391  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[41] ), .O(\edb_top_inst/la0/n1326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4391 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4392  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[42] ), .O(\edb_top_inst/la0/n1327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4392 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4393  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n3180 ), 
            .O(\edb_top_inst/n3183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4393 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4394  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .I3(\edb_top_inst/n3175 ), .O(\edb_top_inst/n3184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4394 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4395  (.I0(\edb_top_inst/n3183 ), .I1(\edb_top_inst/n3184 ), 
            .O(\edb_top_inst/la0/n1381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4395 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4396  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n3180 ), 
            .I3(\edb_top_inst/n3184 ), .O(\edb_top_inst/la0/n1898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4396 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4397  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/edb_user_dr[63] ), 
            .I3(\edb_top_inst/edb_user_dr[66] ), .O(\edb_top_inst/n3185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4397 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4398  (.I0(\edb_top_inst/n3179 ), .I1(\edb_top_inst/n3184 ), 
            .I2(\edb_top_inst/n3185 ), .O(\edb_top_inst/la0/n1950 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4398 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4399  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(\edb_top_inst/la0/address_counter[9] ), .I2(\edb_top_inst/la0/address_counter[10] ), 
            .I3(\edb_top_inst/la0/address_counter[11] ), .O(\edb_top_inst/n3186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4399 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4400  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/la0/address_counter[12] ), .I2(\edb_top_inst/la0/address_counter[13] ), 
            .I3(\edb_top_inst/la0/address_counter[14] ), .O(\edb_top_inst/n3187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4400 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4401  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(\edb_top_inst/la0/address_counter[5] ), .I2(\edb_top_inst/la0/address_counter[6] ), 
            .I3(\edb_top_inst/la0/address_counter[7] ), .O(\edb_top_inst/n3188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4401 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4402  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/address_counter[1] ), .I2(\edb_top_inst/la0/address_counter[2] ), 
            .O(\edb_top_inst/n3189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4402 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4403  (.I0(\edb_top_inst/n3186 ), .I1(\edb_top_inst/n3187 ), 
            .I2(\edb_top_inst/n3188 ), .I3(\edb_top_inst/n3189 ), .O(\edb_top_inst/n3190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4403 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4404  (.I0(\edb_top_inst/n3190 ), .I1(\edb_top_inst/n59 ), 
            .I2(\edb_top_inst/edb_user_dr[45] ), .I3(\edb_top_inst/n3178 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4404 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4405  (.I0(\edb_top_inst/la0/module_next_state[0] ), 
            .I1(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4405 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4406  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[0] ), 
            .I3(\edb_top_inst/la0/biu_ready ), .O(\edb_top_inst/n3191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4406 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4407  (.I0(\edb_top_inst/n3144 ), .I1(\edb_top_inst/n3191 ), 
            .O(\edb_top_inst/n3192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4407 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4408  (.I0(\edb_top_inst/la0/word_count[1] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/la0/word_count[3] ), 
            .O(\edb_top_inst/n3193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4408 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4409  (.I0(\edb_top_inst/n3137 ), .I1(\edb_top_inst/n3138 ), 
            .I2(\edb_top_inst/n3139 ), .I3(\edb_top_inst/n3193 ), .O(\edb_top_inst/n3194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4409 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4410  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n3195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4410 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4411  (.I0(\edb_top_inst/n3192 ), .I1(\edb_top_inst/la0/word_count[0] ), 
            .I2(\edb_top_inst/n3195 ), .I3(\edb_top_inst/n3194 ), .O(\edb_top_inst/n3196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4411 .LUTMASK = 16'h3f05;
    EFX_LUT4 \edb_top_inst/LUT__4412  (.I0(\edb_top_inst/n3151 ), .I1(\edb_top_inst/n3153 ), 
            .I2(\edb_top_inst/n3155 ), .O(\edb_top_inst/n3197 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4412 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4413  (.I0(\edb_top_inst/n3194 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n3198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4413 .LUTMASK = 16'h3001;
    EFX_LUT4 \edb_top_inst/LUT__4414  (.I0(\edb_top_inst/n3198 ), .I1(\edb_top_inst/n3197 ), 
            .I2(\edb_top_inst/n3168 ), .O(\edb_top_inst/n3199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4414 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4415  (.I0(\edb_top_inst/n3196 ), .I1(\edb_top_inst/n3199 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n3200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4415 .LUTMASK = 16'hccca;
    EFX_LUT4 \edb_top_inst/LUT__4416  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3200 ), .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4416 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4417  (.I0(\edb_top_inst/la0/opcode[1] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n1224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4417 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4418  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n3201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4418 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4419  (.I0(\edb_top_inst/n3195 ), .I1(\edb_top_inst/n3146 ), 
            .I2(\edb_top_inst/n3197 ), .I3(\edb_top_inst/n3201 ), .O(\edb_top_inst/n3202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4419 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4420  (.I0(\edb_top_inst/n3170 ), .I1(\edb_top_inst/n3168 ), 
            .I2(\edb_top_inst/n3192 ), .I3(\edb_top_inst/n3202 ), .O(\edb_top_inst/n3203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4420 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__4421  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/n3203 ), .O(\edb_top_inst/la0/n2174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4421 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4422  (.I0(\edb_top_inst/n3146 ), .I1(\edb_top_inst/n3160 ), 
            .I2(\edb_top_inst/n3195 ), .I3(\edb_top_inst/n3201 ), .O(\edb_top_inst/n3204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4422 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__4423  (.I0(\edb_top_inst/n3146 ), .I1(\edb_top_inst/n3173 ), 
            .I2(\edb_top_inst/n3204 ), .I3(\edb_top_inst/n3203 ), .O(\edb_top_inst/ceg_net26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4423 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__4424  (.I0(\edb_top_inst/edb_user_dr[29] ), 
            .I1(\edb_top_inst/la0/word_count[0] ), .I2(\edb_top_inst/n3178 ), 
            .O(\edb_top_inst/la0/data_to_word_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4424 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__4425  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_next_state[0] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/n3203 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4425 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__4426  (.I0(\edb_top_inst/la0/internal_register_select[10] ), 
            .I1(\edb_top_inst/la0/internal_register_select[11] ), .O(\edb_top_inst/n3205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4426 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4427  (.I0(\edb_top_inst/la0/internal_register_select[2] ), 
            .I1(\edb_top_inst/la0/internal_register_select[4] ), .I2(\edb_top_inst/la0/internal_register_select[6] ), 
            .I3(\edb_top_inst/la0/internal_register_select[9] ), .O(\edb_top_inst/n3206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4427 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4428  (.I0(\edb_top_inst/la0/internal_register_select[1] ), 
            .I1(\edb_top_inst/la0/internal_register_select[5] ), .I2(\edb_top_inst/la0/internal_register_select[7] ), 
            .I3(\edb_top_inst/la0/internal_register_select[8] ), .O(\edb_top_inst/n3207 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4428 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4429  (.I0(\edb_top_inst/la0/internal_register_select[12] ), 
            .I1(\edb_top_inst/n3205 ), .I2(\edb_top_inst/n3206 ), .I3(\edb_top_inst/n3207 ), 
            .O(\edb_top_inst/n3208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4429 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4430  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n3209 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec07, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4430 .LUTMASK = 16'hec07;
    EFX_LUT4 \edb_top_inst/LUT__4431  (.I0(\edb_top_inst/n3209 ), .I1(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I2(\edb_top_inst/la0/internal_register_select[3] ), .I3(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4431 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__4432  (.I0(\edb_top_inst/n3161 ), .I1(\edb_top_inst/n3178 ), 
            .O(\edb_top_inst/n3211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4432 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4433  (.I0(\edb_top_inst/n3210 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[1] ), .I3(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4433 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4434  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/n3192 ), .O(\edb_top_inst/n3213 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4434 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4435  (.I0(\edb_top_inst/n3192 ), .I1(\edb_top_inst/n3197 ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .I3(\edb_top_inst/n3213 ), 
            .O(\edb_top_inst/n3214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4435 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__4436  (.I0(\edb_top_inst/n3212 ), .I1(\edb_top_inst/la0/data_from_biu[0] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4436 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4437  (.I0(jtag_inst2_SHIFT), .I1(jtag_inst2_CAPTURE), 
            .I2(\edb_top_inst/n3172 ), .O(\edb_top_inst/n3215 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4437 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4438  (.I0(\edb_top_inst/n3157 ), .I1(\edb_top_inst/n3215 ), 
            .I2(\edb_top_inst/n3213 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/ceg_net14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4438 .LUTMASK = 16'hff70;
    EFX_LUT4 \edb_top_inst/LUT__4439  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/n3181 ), .O(\edb_top_inst/n3216 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4439 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4440  (.I0(\edb_top_inst/n3175 ), .I1(\edb_top_inst/n3216 ), 
            .O(\edb_top_inst/la0/n2751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4440 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4441  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .I3(\edb_top_inst/n3181 ), .O(\edb_top_inst/n3217 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4441 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4442  (.I0(\edb_top_inst/n3175 ), .I1(\edb_top_inst/n3217 ), 
            .O(\edb_top_inst/la0/n3584 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4442 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4443  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n3218 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4443 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4444  (.I0(\edb_top_inst/n3181 ), .I1(\edb_top_inst/n3218 ), 
            .O(\edb_top_inst/n3219 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4444 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4445  (.I0(\edb_top_inst/n3175 ), .I1(\edb_top_inst/n3219 ), 
            .O(\edb_top_inst/la0/n4417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4445 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4446  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n3220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4446 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4447  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/n3220 ), 
            .O(\edb_top_inst/la0/n5250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4447 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4448  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3220 ), 
            .O(\edb_top_inst/la0/n6083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4448 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4449  (.I0(\edb_top_inst/n3217 ), .I1(\edb_top_inst/n3220 ), 
            .O(\edb_top_inst/la0/n6972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4449 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4450  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .I3(\edb_top_inst/n3220 ), .O(\edb_top_inst/n3221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4450 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4451  (.I0(\edb_top_inst/n3183 ), .I1(\edb_top_inst/n3221 ), 
            .O(\edb_top_inst/la0/n6987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4451 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4452  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n3180 ), 
            .O(\edb_top_inst/n3222 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4452 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4453  (.I0(\edb_top_inst/n3221 ), .I1(\edb_top_inst/n3222 ), 
            .O(\edb_top_inst/la0/n7185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4453 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4454  (.I0(\edb_top_inst/n3219 ), .I1(\edb_top_inst/n3220 ), 
            .O(\edb_top_inst/la0/n7869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4454 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4455  (.I0(\edb_top_inst/n3183 ), .I1(\edb_top_inst/n3218 ), 
            .I2(\edb_top_inst/n3220 ), .O(\edb_top_inst/la0/n7884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4455 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4456  (.I0(\edb_top_inst/n3218 ), .I1(\edb_top_inst/n3220 ), 
            .I2(\edb_top_inst/n3222 ), .O(\edb_top_inst/la0/n8082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4456 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4457  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[74] ), .O(\edb_top_inst/n3223 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4457 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4458  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/n3223 ), 
            .O(\edb_top_inst/la0/n8710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4458 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4459  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3223 ), 
            .O(\edb_top_inst/la0/n9543 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4459 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4460  (.I0(\edb_top_inst/n3217 ), .I1(\edb_top_inst/n3223 ), 
            .O(\edb_top_inst/la0/n10376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4460 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4461  (.I0(\edb_top_inst/n3219 ), .I1(\edb_top_inst/n3223 ), 
            .O(\edb_top_inst/la0/n11209 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4461 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4462  (.I0(\edb_top_inst/edb_user_dr[75] ), 
            .I1(\edb_top_inst/edb_user_dr[76] ), .I2(\edb_top_inst/edb_user_dr[73] ), 
            .I3(\edb_top_inst/edb_user_dr[74] ), .O(\edb_top_inst/n3224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4462 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4463  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/n3224 ), 
            .O(\edb_top_inst/la0/n12042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4463 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4464  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3224 ), 
            .O(\edb_top_inst/la0/n12875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4464 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4465  (.I0(\edb_top_inst/n3217 ), .I1(\edb_top_inst/n3224 ), 
            .O(\edb_top_inst/la0/n13708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4465 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4466  (.I0(\edb_top_inst/n3219 ), .I1(\edb_top_inst/n3224 ), 
            .O(\edb_top_inst/la0/n14541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4466 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4467  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[75] ), .O(\edb_top_inst/n3225 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4467 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4468  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3225 ), 
            .O(\edb_top_inst/la0/n16207 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4468 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4469  (.I0(\edb_top_inst/n3217 ), .I1(\edb_top_inst/n3225 ), 
            .O(\edb_top_inst/la0/n17040 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4469 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4470  (.I0(\edb_top_inst/n3219 ), .I1(\edb_top_inst/n3225 ), 
            .O(\edb_top_inst/la0/n17887 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4470 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4471  (.I0(\edb_top_inst/n3183 ), .I1(\edb_top_inst/n3218 ), 
            .I2(\edb_top_inst/n3225 ), .O(\edb_top_inst/la0/n17902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4471 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4472  (.I0(\edb_top_inst/n3218 ), .I1(\edb_top_inst/n3222 ), 
            .I2(\edb_top_inst/n3225 ), .O(\edb_top_inst/la0/n18100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4472 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4473  (.I0(\edb_top_inst/n3167 ), .I1(\edb_top_inst/n3177 ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4473 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4474  (.I0(\edb_top_inst/n3190 ), .I1(\edb_top_inst/n1087 ), 
            .I2(\edb_top_inst/edb_user_dr[46] ), .I3(\edb_top_inst/n3178 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4474 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4475  (.I0(\edb_top_inst/n3190 ), .I1(\edb_top_inst/n1085 ), 
            .I2(\edb_top_inst/edb_user_dr[47] ), .I3(\edb_top_inst/n3178 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4475 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4476  (.I0(\edb_top_inst/n3190 ), .I1(\edb_top_inst/n1083 ), 
            .I2(\edb_top_inst/edb_user_dr[48] ), .I3(\edb_top_inst/n3178 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4476 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4477  (.I0(\edb_top_inst/edb_user_dr[49] ), 
            .I1(\edb_top_inst/n1081 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4477 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4478  (.I0(\edb_top_inst/edb_user_dr[50] ), 
            .I1(\edb_top_inst/n1079 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4478 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4479  (.I0(\edb_top_inst/edb_user_dr[51] ), 
            .I1(\edb_top_inst/n1077 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4479 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4480  (.I0(\edb_top_inst/edb_user_dr[52] ), 
            .I1(\edb_top_inst/n1075 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4480 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4481  (.I0(\edb_top_inst/edb_user_dr[53] ), 
            .I1(\edb_top_inst/n1073 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4481 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4482  (.I0(\edb_top_inst/edb_user_dr[54] ), 
            .I1(\edb_top_inst/n1071 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4482 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4483  (.I0(\edb_top_inst/edb_user_dr[55] ), 
            .I1(\edb_top_inst/n1069 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4483 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4484  (.I0(\edb_top_inst/edb_user_dr[56] ), 
            .I1(\edb_top_inst/n1067 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4484 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4485  (.I0(\edb_top_inst/edb_user_dr[57] ), 
            .I1(\edb_top_inst/n1065 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4485 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4486  (.I0(\edb_top_inst/edb_user_dr[58] ), 
            .I1(\edb_top_inst/n1063 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4486 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4487  (.I0(\edb_top_inst/edb_user_dr[59] ), 
            .I1(\edb_top_inst/n1061 ), .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4487 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4488  (.I0(\edb_top_inst/n1059 ), .I1(\edb_top_inst/la0/address_counter[15] ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3226 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4488 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4489  (.I0(\edb_top_inst/n3226 ), .I1(\edb_top_inst/edb_user_dr[60] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4489 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4490  (.I0(\edb_top_inst/n1202 ), .I1(\edb_top_inst/n1057 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3227 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4490 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4491  (.I0(\edb_top_inst/n3227 ), .I1(\edb_top_inst/edb_user_dr[61] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4491 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4492  (.I0(\edb_top_inst/n1119 ), .I1(\edb_top_inst/n1055 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3228 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4492 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4493  (.I0(\edb_top_inst/n3228 ), .I1(\edb_top_inst/edb_user_dr[62] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4493 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4494  (.I0(\edb_top_inst/n1117 ), .I1(\edb_top_inst/n1053 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3229 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4494 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4495  (.I0(\edb_top_inst/n3229 ), .I1(\edb_top_inst/edb_user_dr[63] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4495 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4496  (.I0(\edb_top_inst/n1115 ), .I1(\edb_top_inst/n1051 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3230 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4496 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4497  (.I0(\edb_top_inst/n3230 ), .I1(\edb_top_inst/edb_user_dr[64] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4497 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4498  (.I0(\edb_top_inst/n1110 ), .I1(\edb_top_inst/n1049 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3231 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4498 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4499  (.I0(\edb_top_inst/n3231 ), .I1(\edb_top_inst/edb_user_dr[65] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4499 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4500  (.I0(\edb_top_inst/n1108 ), .I1(\edb_top_inst/n1047 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3232 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4500 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4501  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/edb_user_dr[66] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4501 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4502  (.I0(\edb_top_inst/n1106 ), .I1(\edb_top_inst/n1045 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4502 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4503  (.I0(\edb_top_inst/n3233 ), .I1(\edb_top_inst/edb_user_dr[67] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4503 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4504  (.I0(\edb_top_inst/n1104 ), .I1(\edb_top_inst/n1043 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4504 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4505  (.I0(\edb_top_inst/n3234 ), .I1(\edb_top_inst/edb_user_dr[68] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4505 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4506  (.I0(\edb_top_inst/n1102 ), .I1(\edb_top_inst/n1041 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3235 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4506 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4507  (.I0(\edb_top_inst/n3235 ), .I1(\edb_top_inst/edb_user_dr[69] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4507 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4508  (.I0(\edb_top_inst/n1100 ), .I1(\edb_top_inst/n1039 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4508 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4509  (.I0(\edb_top_inst/n3236 ), .I1(\edb_top_inst/edb_user_dr[70] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4509 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4510  (.I0(\edb_top_inst/n1098 ), .I1(\edb_top_inst/n1037 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3237 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4510 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4511  (.I0(\edb_top_inst/n3237 ), .I1(\edb_top_inst/edb_user_dr[71] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4511 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4512  (.I0(\edb_top_inst/n1096 ), .I1(\edb_top_inst/n1035 ), 
            .I2(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4512 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4513  (.I0(\edb_top_inst/n3238 ), .I1(\edb_top_inst/edb_user_dr[72] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_addr_counter[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4513 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4522  (.I0(\edb_top_inst/n61 ), .I1(\edb_top_inst/n3203 ), 
            .O(\edb_top_inst/la0/n2173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4522 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4523  (.I0(\edb_top_inst/n1026 ), .I1(\edb_top_inst/n3203 ), 
            .O(\edb_top_inst/la0/n2172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4523 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4524  (.I0(\edb_top_inst/n1024 ), .I1(\edb_top_inst/n3203 ), 
            .O(\edb_top_inst/la0/n2171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4524 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4525  (.I0(\edb_top_inst/n1022 ), .I1(\edb_top_inst/n3203 ), 
            .O(\edb_top_inst/la0/n2170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4525 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4526  (.I0(\edb_top_inst/n1021 ), .I1(\edb_top_inst/n3203 ), 
            .O(\edb_top_inst/la0/n2169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4526 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4527  (.I0(\edb_top_inst/edb_user_dr[30] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[0] ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4527 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__4528  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .O(\edb_top_inst/n3243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4528 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4529  (.I0(\edb_top_inst/edb_user_dr[31] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/n3243 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4529 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4530  (.I0(\edb_top_inst/la0/word_count[2] ), 
            .I1(\edb_top_inst/n3243 ), .I2(\edb_top_inst/la0/word_count[3] ), 
            .O(\edb_top_inst/n3244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4530 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__4531  (.I0(\edb_top_inst/n3244 ), .I1(\edb_top_inst/edb_user_dr[32] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4531 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4532  (.I0(\edb_top_inst/edb_user_dr[33] ), 
            .I1(\edb_top_inst/la0/word_count[4] ), .I2(\edb_top_inst/n3136 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4532 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4533  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/n3136 ), .O(\edb_top_inst/n3245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4533 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4534  (.I0(\edb_top_inst/edb_user_dr[34] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/n3245 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4534 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4535  (.I0(\edb_top_inst/la0/word_count[5] ), 
            .I1(\edb_top_inst/n3245 ), .O(\edb_top_inst/n3246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4535 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4536  (.I0(\edb_top_inst/edb_user_dr[35] ), 
            .I1(\edb_top_inst/la0/word_count[6] ), .I2(\edb_top_inst/n3246 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4536 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4537  (.I0(\edb_top_inst/la0/word_count[6] ), 
            .I1(\edb_top_inst/n3246 ), .O(\edb_top_inst/n3247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4537 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4538  (.I0(\edb_top_inst/edb_user_dr[36] ), 
            .I1(\edb_top_inst/la0/word_count[7] ), .I2(\edb_top_inst/n3247 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4538 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4539  (.I0(\edb_top_inst/n3136 ), .I1(\edb_top_inst/n3137 ), 
            .O(\edb_top_inst/n3248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4539 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4540  (.I0(\edb_top_inst/edb_user_dr[37] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/n3248 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4540 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4541  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/n3248 ), .I2(\edb_top_inst/la0/word_count[9] ), 
            .O(\edb_top_inst/n3249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4541 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__4542  (.I0(\edb_top_inst/n3249 ), .I1(\edb_top_inst/edb_user_dr[38] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4542 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4543  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/la0/word_count[9] ), .I2(\edb_top_inst/n3248 ), 
            .O(\edb_top_inst/n3250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4543 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4544  (.I0(\edb_top_inst/edb_user_dr[39] ), 
            .I1(\edb_top_inst/la0/word_count[10] ), .I2(\edb_top_inst/n3250 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4544 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4545  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/n3250 ), .O(\edb_top_inst/n3251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4545 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4546  (.I0(\edb_top_inst/edb_user_dr[40] ), 
            .I1(\edb_top_inst/la0/word_count[11] ), .I2(\edb_top_inst/n3251 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4546 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4547  (.I0(\edb_top_inst/la0/word_count[11] ), 
            .I1(\edb_top_inst/n3251 ), .O(\edb_top_inst/n3252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4547 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4548  (.I0(\edb_top_inst/edb_user_dr[41] ), 
            .I1(\edb_top_inst/la0/word_count[12] ), .I2(\edb_top_inst/n3252 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4548 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4549  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/la0/word_count[11] ), .I2(\edb_top_inst/la0/word_count[12] ), 
            .I3(\edb_top_inst/n3250 ), .O(\edb_top_inst/n3253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4549 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4550  (.I0(\edb_top_inst/edb_user_dr[42] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/n3253 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4550 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4551  (.I0(\edb_top_inst/n3138 ), .I1(\edb_top_inst/n3250 ), 
            .O(\edb_top_inst/n3254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4551 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4552  (.I0(\edb_top_inst/edb_user_dr[43] ), 
            .I1(\edb_top_inst/la0/word_count[14] ), .I2(\edb_top_inst/n3254 ), 
            .I3(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4552 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4553  (.I0(\edb_top_inst/la0/word_count[14] ), 
            .I1(\edb_top_inst/n3254 ), .I2(\edb_top_inst/la0/word_count[15] ), 
            .O(\edb_top_inst/n3255 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4553 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__4554  (.I0(\edb_top_inst/n3255 ), .I1(\edb_top_inst/edb_user_dr[44] ), 
            .I2(\edb_top_inst/n3178 ), .O(\edb_top_inst/la0/data_to_word_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4554 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4555  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4555 .LUTMASK = 16'hfb8f;
    EFX_LUT4 \edb_top_inst/LUT__4556  (.I0(\edb_top_inst/n3256 ), .I1(\edb_top_inst/la0/la_trig_mask[1] ), 
            .I2(\edb_top_inst/la0/internal_register_select[3] ), .I3(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3257 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4556 .LUTMASK = 16'h030a;
    EFX_LUT4 \edb_top_inst/LUT__4557  (.I0(\edb_top_inst/n3257 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[2] ), .I3(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4557 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4558  (.I0(\edb_top_inst/n3258 ), .I1(\edb_top_inst/la0/data_from_biu[1] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4558 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4559  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n3259 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4559 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4560  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/n3259 ), 
            .O(\edb_top_inst/n3260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4560 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4561  (.I0(\edb_top_inst/n3260 ), .I1(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I2(\edb_top_inst/la0/internal_register_select[3] ), .I3(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3261 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4561 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4562  (.I0(\edb_top_inst/n3261 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[3] ), .I3(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3262 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4562 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4563  (.I0(\edb_top_inst/n3262 ), .I1(\edb_top_inst/la0/data_from_biu[2] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4563 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4564  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/n3208 ), 
            .I3(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3263 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4564 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4565  (.I0(\edb_top_inst/n3208 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4565 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4566  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[3] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4566 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4567  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n3208 ), .O(\edb_top_inst/n3266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4567 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4568  (.I0(\edb_top_inst/n3266 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4568 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4569  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(\edb_top_inst/la0/data_from_biu[3] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4569 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4570  (.I0(\edb_top_inst/n3214 ), .I1(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4570 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4571  (.I0(\edb_top_inst/n3268 ), .I1(\edb_top_inst/n3265 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[4] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4571 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4572  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/data_from_biu[4] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4572 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4573  (.I0(\edb_top_inst/n3208 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/la0/internal_register_select[3] ), .I3(\edb_top_inst/n3214 ), 
            .O(\edb_top_inst/n3271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4573 .LUTMASK = 16'h007d;
    EFX_LUT4 \edb_top_inst/LUT__4574  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[4] ), 
            .I2(\edb_top_inst/n3271 ), .O(\edb_top_inst/n3272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4574 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4575  (.I0(\edb_top_inst/n3272 ), .I1(\edb_top_inst/n3270 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[5] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4575 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4576  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[5] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3266 ), .O(\edb_top_inst/n3273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4576 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4577  (.I0(\edb_top_inst/n3273 ), .I1(\edb_top_inst/la0/data_from_biu[5] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4577 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4578  (.I0(\edb_top_inst/n3274 ), .I1(\edb_top_inst/la0/data_out_shift_reg[6] ), 
            .I2(\edb_top_inst/n3269 ), .O(\edb_top_inst/la0/n2446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4578 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4579  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[6] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4579 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4580  (.I0(\edb_top_inst/n3275 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[7] ), .I3(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4580 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4581  (.I0(\edb_top_inst/n3276 ), .I1(\edb_top_inst/la0/data_from_biu[6] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4581 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4582  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[7] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4582 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4583  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(\edb_top_inst/la0/data_from_biu[7] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4583 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4584  (.I0(\edb_top_inst/n3278 ), .I1(\edb_top_inst/n3277 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[8] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4584 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4585  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3266 ), .O(\edb_top_inst/n3279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4585 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4586  (.I0(\edb_top_inst/n3279 ), .I1(\edb_top_inst/la0/data_from_biu[8] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4586 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4587  (.I0(\edb_top_inst/n3280 ), .I1(\edb_top_inst/la0/data_out_shift_reg[9] ), 
            .I2(\edb_top_inst/n3269 ), .O(\edb_top_inst/la0/n2443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4587 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4588  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[9] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4588 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4589  (.I0(\edb_top_inst/n3281 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[10] ), .I3(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4589 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4590  (.I0(\edb_top_inst/n3282 ), .I1(\edb_top_inst/la0/data_from_biu[9] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4590 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4591  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[10] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3266 ), .O(\edb_top_inst/n3283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4591 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4592  (.I0(\edb_top_inst/n3283 ), .I1(\edb_top_inst/la0/data_from_biu[10] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4592 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4593  (.I0(\edb_top_inst/n3284 ), .I1(\edb_top_inst/la0/data_out_shift_reg[11] ), 
            .I2(\edb_top_inst/n3269 ), .O(\edb_top_inst/la0/n2441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4593 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4594  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[11] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4594 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4595  (.I0(\edb_top_inst/n3285 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[12] ), .I3(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4595 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4596  (.I0(\edb_top_inst/n3286 ), .I1(\edb_top_inst/la0/data_from_biu[11] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4596 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4597  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[12] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4597 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4598  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(\edb_top_inst/la0/data_from_biu[12] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4598 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4599  (.I0(\edb_top_inst/n3288 ), .I1(\edb_top_inst/n3287 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[13] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4599 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4600  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[13] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4600 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4601  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(\edb_top_inst/la0/data_from_biu[13] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4601 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4602  (.I0(\edb_top_inst/n3290 ), .I1(\edb_top_inst/n3289 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[14] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4602 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4603  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(\edb_top_inst/la0/data_from_biu[14] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4603 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4604  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[14] ), 
            .I2(\edb_top_inst/n3271 ), .O(\edb_top_inst/n3292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4604 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4605  (.I0(\edb_top_inst/n3292 ), .I1(\edb_top_inst/n3291 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[15] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4605 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4606  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[15] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4606 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4607  (.I0(\edb_top_inst/la0/la_sample_cnt[12] ), 
            .I1(\edb_top_inst/la0/data_from_biu[15] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4607 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4608  (.I0(\edb_top_inst/n3294 ), .I1(\edb_top_inst/n3293 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[16] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4608 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4609  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[16] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4609 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4610  (.I0(\edb_top_inst/la0/la_sample_cnt[13] ), 
            .I1(\edb_top_inst/la0/data_from_biu[16] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4610 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4611  (.I0(\edb_top_inst/n3296 ), .I1(\edb_top_inst/n3295 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[17] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4611 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4612  (.I0(\edb_top_inst/la0/la_trig_mask[17] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .O(\edb_top_inst/n3297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4612 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4613  (.I0(\edb_top_inst/n3297 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[18] ), .I3(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4613 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4614  (.I0(\edb_top_inst/n3298 ), .I1(\edb_top_inst/la0/data_from_biu[17] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4614 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4615  (.I0(\edb_top_inst/la0/la_trig_mask[18] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .O(\edb_top_inst/n3299 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4615 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4616  (.I0(\edb_top_inst/n3299 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[19] ), .I3(\edb_top_inst/n3211 ), 
            .O(\edb_top_inst/n3300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4616 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4617  (.I0(\edb_top_inst/n3300 ), .I1(\edb_top_inst/la0/data_from_biu[18] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4617 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4618  (.I0(\edb_top_inst/n3211 ), .I1(\edb_top_inst/n3208 ), 
            .O(\edb_top_inst/n3301 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4618 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4619  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/n3301 ), 
            .O(\edb_top_inst/n3302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4619 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4620  (.I0(\edb_top_inst/n3211 ), .I1(\edb_top_inst/la0/data_out_shift_reg[20] ), 
            .I2(\edb_top_inst/la0/data_from_biu[19] ), .I3(\edb_top_inst/n3214 ), 
            .O(\edb_top_inst/n3303 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4620 .LUTMASK = 16'h0fbb;
    EFX_LUT4 \edb_top_inst/LUT__4621  (.I0(\edb_top_inst/la0/la_trig_mask[19] ), 
            .I1(\edb_top_inst/n3302 ), .I2(\edb_top_inst/n3303 ), .O(\edb_top_inst/la0/n2432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4621 .LUTMASK = 16'h8f8f;
    EFX_LUT4 \edb_top_inst/LUT__4622  (.I0(\edb_top_inst/la0/la_trig_mask[20] ), 
            .I1(\edb_top_inst/la0/la_run_trig ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3266 ), .O(\edb_top_inst/n3304 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4622 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4623  (.I0(\edb_top_inst/n3304 ), .I1(\edb_top_inst/la0/data_from_biu[20] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3305 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4623 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4624  (.I0(\edb_top_inst/n3305 ), .I1(\edb_top_inst/la0/data_out_shift_reg[21] ), 
            .I2(\edb_top_inst/n3269 ), .O(\edb_top_inst/la0/n2431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4624 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4625  (.I0(\edb_top_inst/la0/data_from_biu[21] ), 
            .I1(\edb_top_inst/la0/la_run_trig_imdt ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4625 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4626  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[21] ), 
            .I2(\edb_top_inst/n3271 ), .O(\edb_top_inst/n3307 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4626 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4627  (.I0(\edb_top_inst/n3307 ), .I1(\edb_top_inst/n3306 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[22] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4627 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4628  (.I0(\edb_top_inst/la0/data_from_biu[22] ), 
            .I1(\edb_top_inst/la0/la_stop_trig ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3308 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4628 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4629  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[22] ), 
            .I2(\edb_top_inst/n3271 ), .O(\edb_top_inst/n3309 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4629 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4630  (.I0(\edb_top_inst/n3309 ), .I1(\edb_top_inst/n3308 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[23] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4630 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4631  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[23] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4631 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4632  (.I0(\edb_top_inst/la0/data_from_biu[23] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[0] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4632 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4633  (.I0(\edb_top_inst/n3311 ), .I1(\edb_top_inst/n3310 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[24] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4633 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4634  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[24] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4634 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4635  (.I0(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I1(\edb_top_inst/la0/data_from_biu[24] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4635 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4636  (.I0(\edb_top_inst/n3313 ), .I1(\edb_top_inst/n3312 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[25] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4636 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4637  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[25] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3266 ), .O(\edb_top_inst/n3314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4637 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4638  (.I0(\edb_top_inst/n3314 ), .I1(\edb_top_inst/la0/data_from_biu[25] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4638 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4639  (.I0(\edb_top_inst/n3315 ), .I1(\edb_top_inst/la0/data_out_shift_reg[26] ), 
            .I2(\edb_top_inst/n3269 ), .O(\edb_top_inst/la0/n2426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4639 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4640  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/data_from_biu[26] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4640 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4641  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[26] ), 
            .I2(\edb_top_inst/n3271 ), .O(\edb_top_inst/n3317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4641 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4642  (.I0(\edb_top_inst/n3317 ), .I1(\edb_top_inst/n3316 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[27] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4642 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4643  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/data_from_biu[27] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4643 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4644  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[27] ), 
            .I2(\edb_top_inst/n3271 ), .O(\edb_top_inst/n3319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4644 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4645  (.I0(\edb_top_inst/n3319 ), .I1(\edb_top_inst/n3318 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[28] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4645 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4646  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[28] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4646 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4647  (.I0(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I1(\edb_top_inst/la0/data_from_biu[28] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4647 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4648  (.I0(\edb_top_inst/n3321 ), .I1(\edb_top_inst/n3320 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[29] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4648 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4649  (.I0(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[29] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3266 ), .O(\edb_top_inst/n3322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4649 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4650  (.I0(\edb_top_inst/n3322 ), .I1(\edb_top_inst/la0/data_from_biu[29] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4650 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4651  (.I0(\edb_top_inst/n3323 ), .I1(\edb_top_inst/la0/data_out_shift_reg[30] ), 
            .I2(\edb_top_inst/n3269 ), .O(\edb_top_inst/la0/n2422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4651 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4652  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[30] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4652 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4653  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/data_from_biu[30] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4653 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4654  (.I0(\edb_top_inst/n3325 ), .I1(\edb_top_inst/n3324 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[31] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4654 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4655  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[31] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3266 ), .O(\edb_top_inst/n3326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4655 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4656  (.I0(\edb_top_inst/n3326 ), .I1(\edb_top_inst/la0/data_from_biu[31] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4656 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4657  (.I0(\edb_top_inst/n3327 ), .I1(\edb_top_inst/la0/data_out_shift_reg[32] ), 
            .I2(\edb_top_inst/n3269 ), .O(\edb_top_inst/la0/n2420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4657 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4658  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[32] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3266 ), .O(\edb_top_inst/n3328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4658 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4659  (.I0(\edb_top_inst/n3328 ), .I1(\edb_top_inst/la0/data_from_biu[32] ), 
            .I2(\edb_top_inst/n3214 ), .O(\edb_top_inst/n3329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4659 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4660  (.I0(\edb_top_inst/n3329 ), .I1(\edb_top_inst/la0/data_out_shift_reg[33] ), 
            .I2(\edb_top_inst/n3269 ), .O(\edb_top_inst/la0/n2419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4660 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4661  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[33] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4661 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4662  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/la0/data_from_biu[33] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4662 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4663  (.I0(\edb_top_inst/n3331 ), .I1(\edb_top_inst/n3330 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[34] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4663 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4664  (.I0(\edb_top_inst/n3263 ), .I1(\edb_top_inst/la0/la_trig_mask[34] ), 
            .I2(\edb_top_inst/n3264 ), .O(\edb_top_inst/n3332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4664 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4665  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/data_from_biu[34] ), .I2(\edb_top_inst/n3267 ), 
            .I3(\edb_top_inst/n3263 ), .O(\edb_top_inst/n3333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4665 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__4666  (.I0(\edb_top_inst/n3333 ), .I1(\edb_top_inst/n3332 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[35] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4666 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4667  (.I0(\edb_top_inst/n3213 ), .I1(\edb_top_inst/n3208 ), 
            .O(\edb_top_inst/n3334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4667 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4668  (.I0(\edb_top_inst/la0/la_trig_mask[35] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[12] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4668 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__4669  (.I0(\edb_top_inst/n3335 ), .I1(\edb_top_inst/n3334 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[36] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4669 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4670  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[36] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4670 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4671  (.I0(\edb_top_inst/n3336 ), .I1(\edb_top_inst/n3334 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[37] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4671 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4672  (.I0(\edb_top_inst/la0/la_trig_pos[14] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[37] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4672 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4673  (.I0(\edb_top_inst/n3211 ), .I1(\edb_top_inst/la0/data_out_shift_reg[38] ), 
            .O(\edb_top_inst/n3338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4673 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4674  (.I0(\edb_top_inst/n3337 ), .I1(\edb_top_inst/n3301 ), 
            .I2(\edb_top_inst/n3338 ), .I3(\edb_top_inst/n3214 ), .O(\edb_top_inst/la0/n2414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4674 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__4675  (.I0(\edb_top_inst/la0/la_trig_mask[38] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[15] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4675 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__4676  (.I0(\edb_top_inst/n3339 ), .I1(\edb_top_inst/n3334 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[39] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4676 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4677  (.I0(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[39] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4677 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4678  (.I0(\edb_top_inst/n3340 ), .I1(\edb_top_inst/n3334 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[40] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4678 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4679  (.I0(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[40] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4679 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4680  (.I0(\edb_top_inst/n3341 ), .I1(\edb_top_inst/n3301 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[41] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4680 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4681  (.I0(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[41] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n3342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4681 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4682  (.I0(\edb_top_inst/n3342 ), .I1(\edb_top_inst/n3334 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[42] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4682 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4683  (.I0(\edb_top_inst/n3211 ), .I1(\edb_top_inst/n3266 ), 
            .O(\edb_top_inst/n3343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4683 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4684  (.I0(\edb_top_inst/la0/la_trig_mask[42] ), 
            .I1(\edb_top_inst/la0/la_capture_pattern[0] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3343 ), .O(\edb_top_inst/n3344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4684 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4685  (.I0(\edb_top_inst/n3269 ), .I1(\edb_top_inst/la0/data_out_shift_reg[43] ), 
            .I2(\edb_top_inst/n3344 ), .O(\edb_top_inst/la0/n2409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4685 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4686  (.I0(\edb_top_inst/la0/la_capture_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[43] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3343 ), .O(\edb_top_inst/n3345 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4686 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4687  (.I0(\edb_top_inst/n3269 ), .I1(\edb_top_inst/la0/data_out_shift_reg[44] ), 
            .I2(\edb_top_inst/n3345 ), .O(\edb_top_inst/la0/n2408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4687 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4688  (.I0(\edb_top_inst/la0/la_trig_mask[44] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3346 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4688 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__4689  (.I0(\edb_top_inst/n3266 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/n3301 ), .O(\edb_top_inst/n3347 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4689 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4690  (.I0(\edb_top_inst/n3346 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[45] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4690 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4691  (.I0(\edb_top_inst/la0/la_trig_mask[45] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4691 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4692  (.I0(\edb_top_inst/n3348 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[46] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4692 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4693  (.I0(\edb_top_inst/la0/la_trig_mask[46] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3349 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4693 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4694  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n3301 ), .O(\edb_top_inst/n3350 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4694 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4695  (.I0(\edb_top_inst/n3349 ), .I1(\edb_top_inst/n3350 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[47] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4695 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4696  (.I0(\edb_top_inst/la0/la_trig_mask[47] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4696 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4697  (.I0(\edb_top_inst/n3351 ), .I1(\edb_top_inst/n3350 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[48] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4697 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4698  (.I0(\edb_top_inst/la0/la_trig_mask[48] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3352 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4698 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4699  (.I0(\edb_top_inst/n3352 ), .I1(\edb_top_inst/n3350 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[49] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4699 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4700  (.I0(\edb_top_inst/la0/la_trig_mask[49] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3353 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4700 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__4701  (.I0(\edb_top_inst/n3353 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[50] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4701 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4702  (.I0(\edb_top_inst/la0/la_trig_mask[50] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3354 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4702 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4703  (.I0(\edb_top_inst/n3354 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[51] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4703 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4704  (.I0(\edb_top_inst/n3269 ), .I1(\edb_top_inst/la0/data_out_shift_reg[52] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[51] ), .I3(\edb_top_inst/n3302 ), 
            .O(\edb_top_inst/la0/n2400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4704 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__4705  (.I0(\edb_top_inst/la0/la_trig_mask[52] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4705 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4706  (.I0(\edb_top_inst/n3355 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[53] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4706 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4707  (.I0(\edb_top_inst/la0/la_trig_mask[53] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3356 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4707 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__4708  (.I0(\edb_top_inst/n3356 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[54] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4708 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4709  (.I0(\edb_top_inst/la0/la_trig_mask[54] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3357 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4709 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4710  (.I0(\edb_top_inst/n3357 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[55] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2397 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4710 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4711  (.I0(\edb_top_inst/la0/la_trig_mask[55] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4711 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4712  (.I0(\edb_top_inst/n3358 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[56] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4712 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4713  (.I0(\edb_top_inst/la0/la_trig_mask[56] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3359 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4713 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4714  (.I0(\edb_top_inst/n3359 ), .I1(\edb_top_inst/n3350 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[57] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2395 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4714 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4715  (.I0(\edb_top_inst/la0/la_trig_mask[57] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3360 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4715 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__4716  (.I0(\edb_top_inst/n3360 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[58] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4716 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4717  (.I0(\edb_top_inst/n3269 ), .I1(\edb_top_inst/la0/data_out_shift_reg[59] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[58] ), .I3(\edb_top_inst/n3302 ), 
            .O(\edb_top_inst/la0/n2393 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4717 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__4718  (.I0(\edb_top_inst/n3269 ), .I1(\edb_top_inst/la0/data_out_shift_reg[60] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[59] ), .I3(\edb_top_inst/n3302 ), 
            .O(\edb_top_inst/la0/n2392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4718 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__4719  (.I0(\edb_top_inst/la0/la_trig_mask[60] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n3361 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4719 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__4720  (.I0(\edb_top_inst/n3361 ), .I1(\edb_top_inst/n3347 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[61] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2391 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4720 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4721  (.I0(\edb_top_inst/la0/la_trig_mask[61] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3362 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4721 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4722  (.I0(\edb_top_inst/n3362 ), .I1(\edb_top_inst/n3350 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[62] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4722 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4723  (.I0(\edb_top_inst/la0/la_trig_mask[62] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n3363 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4723 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4724  (.I0(\edb_top_inst/n3363 ), .I1(\edb_top_inst/n3350 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[63] ), .I3(\edb_top_inst/n3269 ), 
            .O(\edb_top_inst/la0/n2389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4724 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4725  (.I0(\edb_top_inst/la0/la_trig_mask[63] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n3301 ), .O(\edb_top_inst/la0/n2388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4725 .LUTMASK = 16'h2c00;
    EFX_LUT4 \edb_top_inst/LUT__4726  (.I0(\edb_top_inst/n3195 ), .I1(\edb_top_inst/n3140 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/n3164 ), 
            .O(\edb_top_inst/n3364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4726 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__4727  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(jtag_inst2_UPDATE), .I2(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n3365 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4727 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4728  (.I0(\edb_top_inst/n3140 ), .I1(\edb_top_inst/n3195 ), 
            .I2(\edb_top_inst/n3161 ), .I3(\edb_top_inst/n3365 ), .O(\edb_top_inst/n3366 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4728 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__4729  (.I0(\edb_top_inst/n3195 ), .I1(\edb_top_inst/n3144 ), 
            .O(\edb_top_inst/n3367 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4729 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4730  (.I0(\edb_top_inst/n3366 ), .I1(\edb_top_inst/n3364 ), 
            .I2(\edb_top_inst/n3367 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/la0/module_next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4730 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4731  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/n3197 ), 
            .I3(\edb_top_inst/n3140 ), .O(\edb_top_inst/n3368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4731 .LUTMASK = 16'hb200;
    EFX_LUT4 \edb_top_inst/LUT__4732  (.I0(\edb_top_inst/n3195 ), .I1(jtag_inst2_UPDATE), 
            .I2(\edb_top_inst/n3201 ), .O(\edb_top_inst/n3369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4732 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4733  (.I0(\edb_top_inst/n3140 ), .I1(\edb_top_inst/n3172 ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .I3(\edb_top_inst/n3144 ), 
            .O(\edb_top_inst/n3370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4733 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4734  (.I0(\edb_top_inst/n3369 ), .I1(\edb_top_inst/n3368 ), 
            .I2(\edb_top_inst/n3192 ), .I3(\edb_top_inst/n3370 ), .O(\edb_top_inst/la0/module_next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4734 .LUTMASK = 16'hfff2;
    EFX_LUT4 \edb_top_inst/LUT__4735  (.I0(\edb_top_inst/n3202 ), .I1(\edb_top_inst/n3172 ), 
            .I2(\edb_top_inst/n3140 ), .I3(\edb_top_inst/n3173 ), .O(\edb_top_inst/n3371 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c5f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4735 .LUTMASK = 16'h0c5f;
    EFX_LUT4 \edb_top_inst/LUT__4736  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/n3371 ), 
            .O(\edb_top_inst/la0/module_next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4736 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4737  (.I0(\edb_top_inst/la0/crc_data_out[1] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4737 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4738  (.I0(\edb_top_inst/n3195 ), .I1(\edb_top_inst/n3173 ), 
            .I2(\edb_top_inst/la0/op_reg_en ), .I3(\edb_top_inst/n3204 ), 
            .O(\edb_top_inst/ceg_net221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4738 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4739  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4739 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4740  (.I0(\edb_top_inst/la0/crc_data_out[3] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4740 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4741  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4741 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4742  (.I0(\edb_top_inst/la0/crc_data_out[5] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4742 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4743  (.I0(jtag_inst2_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I2(\edb_top_inst/la0/crc_data_out[0] ), .I3(\edb_top_inst/n3172 ), 
            .O(\edb_top_inst/n3372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3a5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4743 .LUTMASK = 16'hc3a5;
    EFX_LUT4 \edb_top_inst/LUT__4744  (.I0(\edb_top_inst/n3195 ), .I1(\edb_top_inst/n3372 ), 
            .I2(\edb_top_inst/n3201 ), .O(\edb_top_inst/n3373 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4744 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4745  (.I0(\edb_top_inst/n3146 ), .I1(\edb_top_inst/n3160 ), 
            .I2(\edb_top_inst/n3373 ), .O(\edb_top_inst/n3374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4745 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__4746  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[6] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4746 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4747  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4747 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4748  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4748 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4749  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[9] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4749 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4750  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[10] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4750 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4751  (.I0(\edb_top_inst/la0/crc_data_out[11] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4751 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4752  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4752 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4753  (.I0(\edb_top_inst/la0/crc_data_out[13] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4753 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4754  (.I0(\edb_top_inst/la0/crc_data_out[14] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4754 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4755  (.I0(\edb_top_inst/la0/crc_data_out[15] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4755 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4756  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[16] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4756 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4757  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4757 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4758  (.I0(\edb_top_inst/la0/crc_data_out[18] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4758 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4759  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4759 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4760  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[20] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4760 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4761  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[21] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4761 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4762  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[22] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4762 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4763  (.I0(\edb_top_inst/la0/crc_data_out[23] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4763 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4764  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[24] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4764 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4765  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[25] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4765 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4766  (.I0(\edb_top_inst/la0/crc_data_out[26] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4766 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4767  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[27] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4767 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4768  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[28] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4768 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4769  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4769 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4770  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[30] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4770 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4771  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[31] ), .I2(\edb_top_inst/n3374 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4771 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4772  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3374 ), .O(\edb_top_inst/la0/axi_crc_i/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4772 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4773  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4773 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4774  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4774 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4775  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4775 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4776  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4776 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4777  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3375 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4777 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4778  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3375 ), .O(\edb_top_inst/n3376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4778 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4779  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3377 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4779 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4780  (.I0(\edb_top_inst/n3377 ), .I1(\edb_top_inst/n3376 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4780 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4781  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4781 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4782  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4782 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4783  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4783 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4784  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4784 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4785  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3378 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4785 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4786  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3378 ), .O(\edb_top_inst/n3379 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4786 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4787  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4787 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4788  (.I0(\edb_top_inst/n3380 ), .I1(\edb_top_inst/n3379 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4788 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4789  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4789 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4790  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4790 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4791  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4791 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4792  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4792 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4793  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4793 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4794  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3381 ), .O(\edb_top_inst/n3382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4794 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4795  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4795 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4796  (.I0(\edb_top_inst/n3383 ), .I1(\edb_top_inst/n3382 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4796 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4797  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4797 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4798  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4798 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4799  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4799 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4800  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4800 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4801  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4801 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4802  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3384 ), .O(\edb_top_inst/n3385 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4802 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4803  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4803 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4804  (.I0(\edb_top_inst/n3386 ), .I1(\edb_top_inst/n3385 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4804 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4805  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4805 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4806  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4806 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4807  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4807 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4808  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4808 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4809  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4809 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4810  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3387 ), .O(\edb_top_inst/n3388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4810 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4811  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4811 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4812  (.I0(\edb_top_inst/n3389 ), .I1(\edb_top_inst/n3388 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4812 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4813  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4813 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4814  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4814 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4815  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), .O(\edb_top_inst/n3390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4815 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4816  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/n3390 ), .O(\edb_top_inst/n3391 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4816 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4817  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/n3391 ), .O(\edb_top_inst/n3392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4817 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4818  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/n3392 ), .O(\edb_top_inst/n3393 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4818 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4819  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] ), 
            .I1(\edb_top_inst/n3393 ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n3394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4819 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4820  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/n3394 ), .O(\edb_top_inst/n3395 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4820 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4821  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/n3395 ), .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4821 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4822  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n3396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4822 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4823  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/n3397 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4823 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4824  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4824 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4825  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4825 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4826  (.I0(\edb_top_inst/n3396 ), .I1(\edb_top_inst/n3397 ), 
            .I2(\edb_top_inst/n3398 ), .I3(\edb_top_inst/n3399 ), .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4826 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4827  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4827 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4828  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4828 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4829  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4829 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4830  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4830 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4831  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n3404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4831 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4832  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4832 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4833  (.I0(\edb_top_inst/n3402 ), .I1(\edb_top_inst/n3403 ), 
            .I2(\edb_top_inst/n3404 ), .I3(\edb_top_inst/n3405 ), .O(\edb_top_inst/n3406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4833 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4834  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/n3401 ), .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3406 ), .O(\edb_top_inst/n3407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h752f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4834 .LUTMASK = 16'h752f;
    EFX_LUT4 \edb_top_inst/LUT__4835  (.I0(\edb_top_inst/n3407 ), .I1(\edb_top_inst/n3400 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4835 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4836  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4836 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4837  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4837 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4838  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4838 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4839  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4839 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4840  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4840 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4841  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4841 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4842  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4842 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4843  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4843 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4844  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4844 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4845  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4845 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4846  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4846 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4847  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4847 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4848  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4848 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4849  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4849 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4850  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4850 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4851  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4851 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4852  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), .O(\edb_top_inst/n3408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4852 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4853  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/n3408 ), .O(\edb_top_inst/n3409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4853 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4854  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/n3409 ), .O(\edb_top_inst/n3410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4854 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4855  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n3411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4855 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4856  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/n3410 ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/n3411 ), .O(\edb_top_inst/n3412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4856 .LUTMASK = 16'hd400;
    EFX_LUT4 \edb_top_inst/LUT__4857  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n3413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4857 .LUTMASK = 16'h8eaf;
    EFX_LUT4 \edb_top_inst/LUT__4858  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/n3412 ), .I3(\edb_top_inst/n3413 ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b22, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4858 .LUTMASK = 16'h2b22;
    EFX_LUT4 \edb_top_inst/LUT__4859  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/n3414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4859 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4860  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4860 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4861  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4861 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4862  (.I0(\edb_top_inst/n3411 ), .I1(\edb_top_inst/n3414 ), 
            .I2(\edb_top_inst/n3415 ), .I3(\edb_top_inst/n3416 ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4862 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4863  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4863 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4864  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4864 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4865  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4865 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4866  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4866 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4867  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n3421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4867 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4868  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4868 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4869  (.I0(\edb_top_inst/n3419 ), .I1(\edb_top_inst/n3420 ), 
            .I2(\edb_top_inst/n3421 ), .I3(\edb_top_inst/n3422 ), .O(\edb_top_inst/n3423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4869 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4870  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/n3418 ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3423 ), .O(\edb_top_inst/n3424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h752f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4870 .LUTMASK = 16'h752f;
    EFX_LUT4 \edb_top_inst/LUT__4871  (.I0(\edb_top_inst/n3424 ), .I1(\edb_top_inst/n3417 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4871 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4872  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4872 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4873  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4873 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4874  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4874 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4875  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4875 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4876  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4876 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4877  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4877 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4878  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4878 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4879  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4879 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4880  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4880 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4881  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4881 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4882  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4882 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4883  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4883 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4884  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4884 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4885  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4885 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4886  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4886 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4887  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4887 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4888  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4888 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4889  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4889 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4890  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4890 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4891  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3425 ), .O(\edb_top_inst/n3426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4891 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4892  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4892 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4893  (.I0(\edb_top_inst/n3427 ), .I1(\edb_top_inst/n3426 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4893 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4894  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4894 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4895  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4895 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4896  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4896 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4897  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4897 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4898  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4898 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4899  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3428 ), .O(\edb_top_inst/n3429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4899 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4900  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4900 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4901  (.I0(\edb_top_inst/n3430 ), .I1(\edb_top_inst/n3429 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4901 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4902  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4902 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4903  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4903 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4904  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4904 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4905  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4905 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4906  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4906 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4907  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3431 ), .O(\edb_top_inst/n3432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4907 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4908  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4908 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4909  (.I0(\edb_top_inst/n3433 ), .I1(\edb_top_inst/n3432 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4909 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4910  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4910 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4911  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4911 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4912  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4912 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4913  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4913 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4914  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4914 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4915  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3434 ), .O(\edb_top_inst/n3435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4915 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4916  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4916 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4917  (.I0(\edb_top_inst/n3436 ), .I1(\edb_top_inst/n3435 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4917 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4918  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4918 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4919  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4919 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4920  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4920 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4921  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4921 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4922  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4922 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4923  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3437 ), .O(\edb_top_inst/n3438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4923 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4924  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4924 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4925  (.I0(\edb_top_inst/n3439 ), .I1(\edb_top_inst/n3438 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4925 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4926  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4926 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4927  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4927 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4928  (.I0(\edb_top_inst/la0/GEN_PROBE[12].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4928 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4929  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4929 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4930  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4930 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4931  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3440 ), .O(\edb_top_inst/n3441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4931 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4932  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4932 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4933  (.I0(\edb_top_inst/n3442 ), .I1(\edb_top_inst/n3441 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[12].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4933 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4934  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4934 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4935  (.I0(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4935 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4936  (.I0(\edb_top_inst/la0/GEN_PROBE[13].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4936 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4937  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4937 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4938  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4938 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4939  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3443 ), .O(\edb_top_inst/n3444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4939 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4940  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4940 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4941  (.I0(\edb_top_inst/n3445 ), .I1(\edb_top_inst/n3444 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[13].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4941 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4942  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4942 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4943  (.I0(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4943 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4944  (.I0(\edb_top_inst/la0/GEN_PROBE[14].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4944 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4945  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4945 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4946  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4946 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4947  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3446 ), .O(\edb_top_inst/n3447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4947 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4948  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4948 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4949  (.I0(\edb_top_inst/n3448 ), .I1(\edb_top_inst/n3447 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[14].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4949 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4950  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/n3225 ), 
            .O(\edb_top_inst/la0/n15374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4950 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4951  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4951 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4952  (.I0(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4952 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4953  (.I0(\edb_top_inst/la0/GEN_PROBE[15].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4953 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4954  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4954 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4955  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4955 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4956  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3449 ), .O(\edb_top_inst/n3450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4956 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4957  (.I0(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4957 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4958  (.I0(\edb_top_inst/n3451 ), .I1(\edb_top_inst/n3450 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[15].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4958 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4959  (.I0(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4959 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4960  (.I0(\edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4960 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4961  (.I0(\edb_top_inst/la0/GEN_PROBE[16].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4961 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4962  (.I0(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4962 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4963  (.I0(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4963 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4964  (.I0(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3452 ), .O(\edb_top_inst/n3453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4964 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4965  (.I0(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4965 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4966  (.I0(\edb_top_inst/n3454 ), .I1(\edb_top_inst/n3453 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[16].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4966 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4967  (.I0(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4967 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4968  (.I0(\edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4968 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4969  (.I0(\edb_top_inst/la0/GEN_PROBE[17].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4969 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4970  (.I0(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4970 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4971  (.I0(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4971 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__4972  (.I0(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n3455 ), .O(\edb_top_inst/n3456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4972 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4973  (.I0(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4973 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__4974  (.I0(\edb_top_inst/n3457 ), .I1(\edb_top_inst/n3456 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[17].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4974 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4975  (.I0(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4975 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4976  (.I0(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4976 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4977  (.I0(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b22, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4977 .LUTMASK = 16'h2b22;
    EFX_LUT4 \edb_top_inst/LUT__4978  (.I0(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/equal_9/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ff6, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4978 .LUTMASK = 16'h6ff6;
    EFX_LUT4 \edb_top_inst/LUT__4979  (.I0(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4979 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4980  (.I0(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n3458 ), .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4980 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4981  (.I0(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4981 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4982  (.I0(\edb_top_inst/n3458 ), .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3460 ), .O(\edb_top_inst/n3461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4c70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4982 .LUTMASK = 16'h4c70;
    EFX_LUT4 \edb_top_inst/LUT__4983  (.I0(\edb_top_inst/n3461 ), .I1(\edb_top_inst/n3459 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4983 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4984  (.I0(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4984 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4985  (.I0(\edb_top_inst/la0/GEN_PROBE[18].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.trigger_cu/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4985 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4986  (.I0(\edb_top_inst/la0/la_trig_mask[18] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[4] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4986 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4987  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[13] ), .I2(\edb_top_inst/n3462 ), 
            .O(\edb_top_inst/n3463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4987 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__4988  (.I0(\edb_top_inst/la0/la_trig_mask[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4988 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4989  (.I0(\edb_top_inst/la0/la_trig_mask[16] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[12] ), .I3(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4989 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4990  (.I0(\edb_top_inst/la0/la_trig_mask[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4990 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4991  (.I0(\edb_top_inst/la0/la_trig_mask[17] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4991 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4992  (.I0(\edb_top_inst/n3464 ), .I1(\edb_top_inst/n3465 ), 
            .I2(\edb_top_inst/n3466 ), .I3(\edb_top_inst/n3467 ), .O(\edb_top_inst/n3468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4992 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4993  (.I0(\edb_top_inst/la0/la_trig_mask[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[10] ), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4993 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4994  (.I0(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4994 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4995  (.I0(\edb_top_inst/la0/la_trig_mask[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4995 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4996  (.I0(\edb_top_inst/la0/la_trig_mask[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4996 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4997  (.I0(\edb_top_inst/n3469 ), .I1(\edb_top_inst/n3470 ), 
            .I2(\edb_top_inst/n3471 ), .I3(\edb_top_inst/n3472 ), .O(\edb_top_inst/n3473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4997 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4998  (.I0(\edb_top_inst/n3463 ), .I1(\edb_top_inst/n3468 ), 
            .I2(\edb_top_inst/n3473 ), .O(\edb_top_inst/n3474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4998 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4999  (.I0(\edb_top_inst/la0/GEN_PROBE[16].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[16] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[3] ), .O(\edb_top_inst/n3475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4999 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5000  (.I0(\edb_top_inst/la0/GEN_PROBE[12].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[12] ), .I2(\edb_top_inst/n3475 ), 
            .O(\edb_top_inst/n3476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5000 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__5001  (.I0(\edb_top_inst/la0/GEN_PROBE[17].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[17] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[4] ), .O(\edb_top_inst/n3477 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5001 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5002  (.I0(\edb_top_inst/la0/GEN_PROBE[18].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[18] ), .I2(\edb_top_inst/la0/GEN_PROBE[15].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[15] ), .O(\edb_top_inst/n3478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5002 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5003  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[8] ), .O(\edb_top_inst/n3479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5003 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5004  (.I0(\edb_top_inst/la0/GEN_PROBE[13].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[9] ), .O(\edb_top_inst/n3480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5004 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5005  (.I0(\edb_top_inst/n3477 ), .I1(\edb_top_inst/n3478 ), 
            .I2(\edb_top_inst/n3479 ), .I3(\edb_top_inst/n3480 ), .O(\edb_top_inst/n3481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5005 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5006  (.I0(\edb_top_inst/la0/GEN_PROBE[14].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[14] ), .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[7] ), .O(\edb_top_inst/n3482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5006 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5007  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[2] ), .O(\edb_top_inst/n3483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5007 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5008  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[10] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[1] ), .O(\edb_top_inst/n3484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5008 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5009  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[6] ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[0] ), .O(\edb_top_inst/n3485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5009 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__5010  (.I0(\edb_top_inst/n3482 ), .I1(\edb_top_inst/n3483 ), 
            .I2(\edb_top_inst/n3484 ), .I3(\edb_top_inst/n3485 ), .O(\edb_top_inst/n3486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5010 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5011  (.I0(\edb_top_inst/n3476 ), .I1(\edb_top_inst/n3481 ), 
            .I2(\edb_top_inst/n3486 ), .O(\edb_top_inst/n3487 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5011 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5012  (.I0(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .I1(\edb_top_inst/n3474 ), .I2(\edb_top_inst/n3487 ), .I3(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .O(\edb_top_inst/la0/trigger_tu/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d32, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5012 .LUTMASK = 16'h0d32;
    EFX_LUT4 \edb_top_inst/LUT__5013  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5013 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5014  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/n3488 ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[12] ), .O(\edb_top_inst/n3489 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfc8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5014 .LUTMASK = 16'hbfc8;
    EFX_LUT4 \edb_top_inst/LUT__5015  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5015 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__5016  (.I0(\edb_top_inst/n3490 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[12] ), 
            .O(\edb_top_inst/n3491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5016 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5017  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3489 ), .I2(\edb_top_inst/n3491 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13] ), 
            .O(\edb_top_inst/n3492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5017 .LUTMASK = 16'h0fee;
    EFX_LUT4 \edb_top_inst/LUT__5018  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5018 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5019  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3493 ), .I2(\edb_top_inst/n3488 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .O(\edb_top_inst/n3494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h45fe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5019 .LUTMASK = 16'h45fe;
    EFX_LUT4 \edb_top_inst/LUT__5020  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5020 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5021  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5021 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5022  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I1(\edb_top_inst/n3495 ), .I2(\edb_top_inst/n3496 ), .O(\edb_top_inst/n3497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5022 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5023  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5023 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5024  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5024 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5025  (.I0(\edb_top_inst/n3498 ), .I1(\edb_top_inst/n3499 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), .O(\edb_top_inst/n3500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5025 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__5026  (.I0(\edb_top_inst/n3497 ), .I1(\edb_top_inst/n3494 ), 
            .I2(\edb_top_inst/n3500 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .O(\edb_top_inst/n3501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5026 .LUTMASK = 16'h030a;
    EFX_LUT4 \edb_top_inst/LUT__5027  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5027 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__5028  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(\edb_top_inst/n3502 ), .O(\edb_top_inst/n3503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5028 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5029  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5029 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5030  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3504 ), .I2(\edb_top_inst/n3495 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n3505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd02f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5030 .LUTMASK = 16'hd02f;
    EFX_LUT4 \edb_top_inst/LUT__5031  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5031 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5032  (.I0(\edb_top_inst/n3506 ), .I1(\edb_top_inst/n3495 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), .O(\edb_top_inst/n3507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5032 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__5033  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5033 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__5034  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .I2(\edb_top_inst/n3508 ), 
            .I3(\edb_top_inst/n3499 ), .O(\edb_top_inst/n3509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5034 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__5035  (.I0(\edb_top_inst/n3503 ), .I1(\edb_top_inst/n3505 ), 
            .I2(\edb_top_inst/n3507 ), .I3(\edb_top_inst/n3509 ), .O(\edb_top_inst/n3510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5035 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__5036  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5036 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5037  (.I0(\edb_top_inst/n3511 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .I3(\edb_top_inst/n3495 ), 
            .O(\edb_top_inst/n3512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5037 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__5038  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n3511 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .O(\edb_top_inst/n3513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf20d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5038 .LUTMASK = 16'hf20d;
    EFX_LUT4 \edb_top_inst/LUT__5039  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5039 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__5040  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3514 ), .O(\edb_top_inst/n3515 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5040 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5041  (.I0(\edb_top_inst/n3512 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I2(\edb_top_inst/n3515 ), .I3(\edb_top_inst/n3513 ), .O(\edb_top_inst/n3516 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5041 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__5042  (.I0(\edb_top_inst/n3492 ), .I1(\edb_top_inst/n3501 ), 
            .I2(\edb_top_inst/n3510 ), .I3(\edb_top_inst/n3516 ), .O(\edb_top_inst/n3517 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5042 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5043  (.I0(\edb_top_inst/n3506 ), .I1(\edb_top_inst/n3495 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n3518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5043 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__5044  (.I0(\edb_top_inst/n3496 ), .I1(\edb_top_inst/n3495 ), 
            .I2(\edb_top_inst/n3518 ), .I3(\edb_top_inst/la0/la_trig_pos[1] ), 
            .O(\edb_top_inst/n3519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5044 .LUTMASK = 16'h0708;
    EFX_LUT4 \edb_top_inst/LUT__5045  (.I0(\edb_top_inst/n3493 ), .I1(\edb_top_inst/n3514 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n3520 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5045 .LUTMASK = 16'h53fc;
    EFX_LUT4 \edb_top_inst/LUT__5046  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3504 ), .I2(\edb_top_inst/n3495 ), .I3(\edb_top_inst/la0/la_trig_pos[4] ), 
            .O(\edb_top_inst/n3521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd02f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5046 .LUTMASK = 16'hd02f;
    EFX_LUT4 \edb_top_inst/LUT__5047  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[16] ), .I2(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3522 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ffc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5047 .LUTMASK = 16'h6ffc;
    EFX_LUT4 \edb_top_inst/LUT__5048  (.I0(\edb_top_inst/n3520 ), .I1(\edb_top_inst/n3521 ), 
            .I2(\edb_top_inst/n3522 ), .O(\edb_top_inst/n3523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5048 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5049  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[7] ), .I2(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I3(\edb_top_inst/n3495 ), .O(\edb_top_inst/n3524 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5049 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__5050  (.I0(\edb_top_inst/n3504 ), .I1(\edb_top_inst/n3488 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[12] ), 
            .O(\edb_top_inst/n3525 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5050 .LUTMASK = 16'hf40b;
    EFX_LUT4 \edb_top_inst/LUT__5051  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/n3502 ), .O(\edb_top_inst/n3526 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5051 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5052  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/n3490 ), .O(\edb_top_inst/n3527 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5052 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5053  (.I0(\edb_top_inst/n3524 ), .I1(\edb_top_inst/n3526 ), 
            .I2(\edb_top_inst/n3527 ), .I3(\edb_top_inst/n3525 ), .O(\edb_top_inst/n3528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5053 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__5054  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5054 .LUTMASK = 16'h7ff8;
    EFX_LUT4 \edb_top_inst/LUT__5055  (.I0(\edb_top_inst/n3498 ), .I1(\edb_top_inst/n3529 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[2] ), .O(\edb_top_inst/n3530 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5055 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__5056  (.I0(\edb_top_inst/n3499 ), .I1(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[14] ), .I3(\edb_top_inst/n3530 ), 
            .O(\edb_top_inst/n3531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbff1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5056 .LUTMASK = 16'hbff1;
    EFX_LUT4 \edb_top_inst/LUT__5057  (.I0(\edb_top_inst/n3531 ), .I1(\edb_top_inst/n3523 ), 
            .I2(\edb_top_inst/n3528 ), .I3(\edb_top_inst/n3519 ), .O(\edb_top_inst/n3532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5057 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5058  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5058 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__5059  (.I0(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[11] ), .I2(\edb_top_inst/n3533 ), 
            .I3(\edb_top_inst/n3508 ), .O(\edb_top_inst/n3534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5059 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__5060  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n3511 ), .O(\edb_top_inst/n3535 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5060 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5061  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/n3511 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[8] ), .O(\edb_top_inst/n3536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe41, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5061 .LUTMASK = 16'hbe41;
    EFX_LUT4 \edb_top_inst/LUT__5062  (.I0(\edb_top_inst/n3535 ), .I1(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[0] ), .I3(\edb_top_inst/n3536 ), 
            .O(\edb_top_inst/n3537 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5062 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__5063  (.I0(\edb_top_inst/n3517 ), .I1(\edb_top_inst/n3532 ), 
            .I2(\edb_top_inst/n3534 ), .I3(\edb_top_inst/n3537 ), .O(\edb_top_inst/n3538 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5063 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5064  (.I0(\edb_top_inst/n3511 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3539 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5064 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__5065  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3514 ), .I2(\edb_top_inst/n3535 ), .O(\edb_top_inst/n3540 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5065 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5066  (.I0(\edb_top_inst/n3539 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .I3(\edb_top_inst/n3540 ), 
            .O(\edb_top_inst/n3541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5066 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__5067  (.I0(\edb_top_inst/n3506 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), .I3(\edb_top_inst/n3495 ), 
            .O(\edb_top_inst/n3542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ecf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5067 .LUTMASK = 16'h1ecf;
    EFX_LUT4 \edb_top_inst/LUT__5068  (.I0(\edb_top_inst/n3511 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I3(\edb_top_inst/n3495 ), 
            .O(\edb_top_inst/n3543 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ecf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5068 .LUTMASK = 16'h7ecf;
    EFX_LUT4 \edb_top_inst/LUT__5069  (.I0(\edb_top_inst/n3542 ), .I1(\edb_top_inst/n3543 ), 
            .O(\edb_top_inst/n3544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5069 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5070  (.I0(\edb_top_inst/n3504 ), .I1(\edb_top_inst/n3499 ), 
            .O(\edb_top_inst/n3545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5070 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5071  (.I0(\edb_top_inst/n3495 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n3504 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n3546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h827f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5071 .LUTMASK = 16'h827f;
    EFX_LUT4 \edb_top_inst/LUT__5072  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(\edb_top_inst/n3545 ), .I2(\edb_top_inst/n3546 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .O(\edb_top_inst/n3547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5072 .LUTMASK = 16'hf0bb;
    EFX_LUT4 \edb_top_inst/LUT__5073  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3548 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5073 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5074  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n3548 ), .O(\edb_top_inst/n3549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5074 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5075  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/n3504 ), .O(\edb_top_inst/n3550 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5415, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5075 .LUTMASK = 16'h5415;
    EFX_LUT4 \edb_top_inst/LUT__5076  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[12] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13] ), 
            .I2(\edb_top_inst/n3549 ), .I3(\edb_top_inst/n3550 ), .O(\edb_top_inst/n3551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5076 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__5077  (.I0(\edb_top_inst/n3511 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/n3533 ), .O(\edb_top_inst/n3552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5077 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__5078  (.I0(\edb_top_inst/n3502 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), .I3(\edb_top_inst/n3552 ), 
            .O(\edb_top_inst/n3553 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5078 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__5079  (.I0(\edb_top_inst/n3499 ), .I1(\edb_top_inst/la0/la_window_depth[0] ), 
            .I2(\edb_top_inst/la0/la_window_depth[1] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .O(\edb_top_inst/n3554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h28d7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5079 .LUTMASK = 16'h28d7;
    EFX_LUT4 \edb_top_inst/LUT__5080  (.I0(\edb_top_inst/n3547 ), .I1(\edb_top_inst/n3551 ), 
            .I2(\edb_top_inst/n3553 ), .I3(\edb_top_inst/n3554 ), .O(\edb_top_inst/n3555 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5080 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5081  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .I2(\edb_top_inst/n3496 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .O(\edb_top_inst/n3556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h30df, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5081 .LUTMASK = 16'h30df;
    EFX_LUT4 \edb_top_inst/LUT__5082  (.I0(\edb_top_inst/n3511 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I2(\edb_top_inst/n3556 ), .I3(\edb_top_inst/n3508 ), .O(\edb_top_inst/n3557 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5082 .LUTMASK = 16'h0b0c;
    EFX_LUT4 \edb_top_inst/LUT__5083  (.I0(\edb_top_inst/n3541 ), .I1(\edb_top_inst/n3544 ), 
            .I2(\edb_top_inst/n3555 ), .I3(\edb_top_inst/n3557 ), .O(\edb_top_inst/n3558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5083 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5084  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[3] ), .O(\edb_top_inst/n3559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5084 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5085  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/la0/la_num_trigger[6] ), 
            .O(\edb_top_inst/n3560 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5085 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5086  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .I2(\edb_top_inst/n3559 ), 
            .I3(\edb_top_inst/n3560 ), .O(\edb_top_inst/n3561 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5086 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5087  (.I0(\edb_top_inst/la0/la_num_trigger[9] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[10] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I3(\edb_top_inst/n3561 ), .O(\edb_top_inst/n3562 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5087 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5088  (.I0(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[9] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I3(\edb_top_inst/n3561 ), .O(\edb_top_inst/n3563 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd33c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5088 .LUTMASK = 16'hd33c;
    EFX_LUT4 \edb_top_inst/LUT__5089  (.I0(\edb_top_inst/n3562 ), .I1(\edb_top_inst/n3563 ), 
            .I2(\edb_top_inst/la0/la_num_trigger[11] ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .O(\edb_top_inst/n3564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc55c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5089 .LUTMASK = 16'hc55c;
    EFX_LUT4 \edb_top_inst/LUT__5090  (.I0(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .O(\edb_top_inst/n3565 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5090 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5091  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .O(\edb_top_inst/n3566 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5091 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5092  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/n3566 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I3(\edb_top_inst/n3559 ), .O(\edb_top_inst/n3567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5092 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__5093  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/n3567 ), 
            .I3(\edb_top_inst/n3565 ), .O(\edb_top_inst/n3568 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b04, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5093 .LUTMASK = 16'h0b04;
    EFX_LUT4 \edb_top_inst/LUT__5094  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[10] ), .O(\edb_top_inst/n3569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5094 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5095  (.I0(\edb_top_inst/la0/la_num_trigger[11] ), 
            .I1(\edb_top_inst/n3559 ), .I2(\edb_top_inst/n3560 ), .I3(\edb_top_inst/n3569 ), 
            .O(\edb_top_inst/n3570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5095 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__5096  (.I0(\edb_top_inst/la0/la_num_trigger[12] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[13] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12] ), 
            .I3(\edb_top_inst/n3570 ), .O(\edb_top_inst/n3571 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5096 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__5097  (.I0(\edb_top_inst/la0/la_num_trigger[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .O(\edb_top_inst/n3572 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5097 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5098  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .O(\edb_top_inst/n3573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5098 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5099  (.I0(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I1(\edb_top_inst/n3572 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I3(\edb_top_inst/n3573 ), .O(\edb_top_inst/n3574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5099 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__5100  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .O(\edb_top_inst/n3575 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5100 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5101  (.I0(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), .O(\edb_top_inst/n3576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5101 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5102  (.I0(\edb_top_inst/n3559 ), .I1(\edb_top_inst/n3560 ), 
            .I2(\edb_top_inst/n3575 ), .I3(\edb_top_inst/n3576 ), .O(\edb_top_inst/n3577 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5102 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__5103  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .O(\edb_top_inst/n3578 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5103 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__5104  (.I0(\edb_top_inst/la0/la_num_trigger[14] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[15] ), .I2(\edb_top_inst/la0/la_num_trigger[16] ), 
            .I3(\edb_top_inst/n3578 ), .O(\edb_top_inst/n3579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5104 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5105  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .O(\edb_top_inst/n3580 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5105 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__5106  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .I2(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .O(\edb_top_inst/n3581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5106 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5107  (.I0(\edb_top_inst/n3580 ), .I1(\edb_top_inst/n3581 ), 
            .I2(\edb_top_inst/n3559 ), .I3(\edb_top_inst/n3560 ), .O(\edb_top_inst/n3582 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha333, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5107 .LUTMASK = 16'ha333;
    EFX_LUT4 \edb_top_inst/LUT__5108  (.I0(\edb_top_inst/n3574 ), .I1(\edb_top_inst/n3582 ), 
            .I2(\edb_top_inst/n3579 ), .I3(\edb_top_inst/n3577 ), .O(\edb_top_inst/n3583 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5108 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5109  (.I0(\edb_top_inst/n3571 ), .I1(\edb_top_inst/n3568 ), 
            .I2(\edb_top_inst/n3583 ), .O(\edb_top_inst/n3584 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5109 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5110  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .I2(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n3585 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5110 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__5111  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[6] ), 
            .O(\edb_top_inst/n3586 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5111 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5112  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[11] ), .O(\edb_top_inst/n3587 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5112 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5113  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .I2(\edb_top_inst/la0/la_trig_pos[9] ), 
            .O(\edb_top_inst/n3588 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5113 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5114  (.I0(\edb_top_inst/n3585 ), .I1(\edb_top_inst/n3586 ), 
            .I2(\edb_top_inst/n3587 ), .I3(\edb_top_inst/n3588 ), .O(\edb_top_inst/n3589 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5114 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5115  (.I0(\edb_top_inst/la0/la_trig_pos[14] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[15] ), .I2(\edb_top_inst/la0/la_trig_pos[16] ), 
            .O(\edb_top_inst/n3590 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5115 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__5116  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[13] ), .I2(\edb_top_inst/n3589 ), 
            .I3(\edb_top_inst/n3590 ), .O(\edb_top_inst/n3591 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5116 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5117  (.I0(\edb_top_inst/n3584 ), .I1(\edb_top_inst/n3564 ), 
            .I2(\edb_top_inst/n3591 ), .O(\edb_top_inst/n3592 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5117 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__5118  (.I0(\edb_top_inst/n3558 ), .I1(\edb_top_inst/n3538 ), 
            .I2(\edb_top_inst/n3592 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3593 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5118 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__5119  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n3594 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5119 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5120  (.I0(\edb_top_inst/n3535 ), .I1(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[0] ), .I3(\edb_top_inst/n3539 ), 
            .O(\edb_top_inst/n3595 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5120 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__5121  (.I0(\edb_top_inst/n3595 ), .I1(\edb_top_inst/n3534 ), 
            .I2(\edb_top_inst/n3532 ), .O(\edb_top_inst/n3596 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5121 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5122  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/la0/la_stop_trig ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n3597 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5122 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__5123  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/n3596 ), 
            .I2(\edb_top_inst/n3597 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3598 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5123 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__5124  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n3599 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5124 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5125  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[9] ), .O(\edb_top_inst/n3600 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5125 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5126  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/n3585 ), .I2(\edb_top_inst/n3586 ), .O(\edb_top_inst/n3601 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5126 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5127  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/n3600 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I3(\edb_top_inst/n3601 ), .O(\edb_top_inst/n3602 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5127 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__5128  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[11] ), .O(\edb_top_inst/n3603 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5128 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5129  (.I0(\edb_top_inst/n3585 ), .I1(\edb_top_inst/n3586 ), 
            .I2(\edb_top_inst/n3588 ), .O(\edb_top_inst/n3604 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5129 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__5130  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/n3603 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I3(\edb_top_inst/n3604 ), .O(\edb_top_inst/n3605 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5130 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__5131  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[12] ), .I2(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I3(\edb_top_inst/n3589 ), .O(\edb_top_inst/n3606 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5131 .LUTMASK = 16'hbac3;
    EFX_LUT4 \edb_top_inst/LUT__5132  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n3607 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5132 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5133  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/n3607 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I3(\edb_top_inst/n3585 ), .O(\edb_top_inst/n3608 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5133 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__5134  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n3609 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5134 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__5135  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n3610 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5135 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5136  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/n3609 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I3(\edb_top_inst/n3610 ), .O(\edb_top_inst/n3611 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5136 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__5137  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I2(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n3612 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5137 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__5138  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n3613 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5138 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__5139  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n3614 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5139 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5140  (.I0(\edb_top_inst/n3612 ), .I1(\edb_top_inst/n3613 ), 
            .I2(\edb_top_inst/n3585 ), .I3(\edb_top_inst/n3614 ), .O(\edb_top_inst/n3615 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha333, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5140 .LUTMASK = 16'ha333;
    EFX_LUT4 \edb_top_inst/LUT__5141  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .O(\edb_top_inst/n3616 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5141 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__5142  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[12] ), .I2(\edb_top_inst/la0/la_trig_pos[13] ), 
            .O(\edb_top_inst/n3617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5142 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__5143  (.I0(\edb_top_inst/n3616 ), .I1(\edb_top_inst/n3617 ), 
            .I2(\edb_top_inst/n3590 ), .O(\edb_top_inst/n3618 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5143 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5144  (.I0(\edb_top_inst/n3608 ), .I1(\edb_top_inst/n3611 ), 
            .I2(\edb_top_inst/n3615 ), .I3(\edb_top_inst/n3618 ), .O(\edb_top_inst/n3619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5144 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__5145  (.I0(\edb_top_inst/n3602 ), .I1(\edb_top_inst/n3605 ), 
            .I2(\edb_top_inst/n3606 ), .I3(\edb_top_inst/n3619 ), .O(\edb_top_inst/n3620 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5145 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5146  (.I0(\edb_top_inst/n3591 ), .I1(\edb_top_inst/n3599 ), 
            .I2(\edb_top_inst/n3620 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3621 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5146 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__5147  (.I0(\edb_top_inst/n3621 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n3622 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5147 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__5148  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n3623 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5148 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__5149  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n3517 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/n3623 ), .O(\edb_top_inst/n3624 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5149 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__5150  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3625 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5150 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5151  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n3626 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5151 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5152  (.I0(\edb_top_inst/n3620 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3626 ), .O(\edb_top_inst/n3627 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5152 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__5153  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3625 ), .I2(\edb_top_inst/n3624 ), .I3(\edb_top_inst/n3627 ), 
            .O(\edb_top_inst/n3628 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5153 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__5154  (.I0(\edb_top_inst/n3593 ), .I1(\edb_top_inst/n3598 ), 
            .I2(\edb_top_inst/n3622 ), .I3(\edb_top_inst/n3628 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5154 .LUTMASK = 16'hb0ff;
    EFX_LUT4 \edb_top_inst/LUT__5155  (.I0(\edb_top_inst/n3200 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/la0/la_biu_inst/n374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5155 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5156  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/n1303 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5156 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5157  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), 
            .I3(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5157 .LUTMASK = 16'h00be;
    EFX_LUT4 \edb_top_inst/LUT__5158  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(\edb_top_inst/ceg_net351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5158 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5159  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/n3596 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3629 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5159 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__5160  (.I0(\edb_top_inst/n3564 ), .I1(\edb_top_inst/n3584 ), 
            .O(\edb_top_inst/n3630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5160 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5161  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3631 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5161 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5162  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3517 ), .O(\edb_top_inst/n3632 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5162 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5163  (.I0(\edb_top_inst/n3630 ), .I1(\edb_top_inst/n3631 ), 
            .I2(\edb_top_inst/n3632 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3633 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5163 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__5164  (.I0(\edb_top_inst/n3593 ), .I1(\edb_top_inst/n3629 ), 
            .I2(\edb_top_inst/n3633 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f44, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5164 .LUTMASK = 16'h0f44;
    EFX_LUT4 \edb_top_inst/LUT__5165  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/n25424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5165 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5166  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/la0/la_stop_trig ), 
            .I2(\edb_top_inst/n3259 ), .O(\edb_top_inst/n3634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5166 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__5167  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/n3596 ), 
            .I2(\edb_top_inst/n3630 ), .I3(\edb_top_inst/n3634 ), .O(\edb_top_inst/n3635 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5167 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__5168  (.I0(\edb_top_inst/n3558 ), .I1(\edb_top_inst/n3538 ), 
            .I2(\edb_top_inst/n3592 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3636 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5168 .LUTMASK = 16'hf100;
    EFX_LUT4 \edb_top_inst/LUT__5169  (.I0(\edb_top_inst/n3256 ), .I1(\edb_top_inst/n3625 ), 
            .O(\edb_top_inst/n3637 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5169 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__5170  (.I0(\edb_top_inst/n3564 ), .I1(\edb_top_inst/n3584 ), 
            .I2(\edb_top_inst/n3631 ), .O(\edb_top_inst/n3638 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5170 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5171  (.I0(\edb_top_inst/n3632 ), .I1(\edb_top_inst/n3638 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I3(\edb_top_inst/n3625 ), 
            .O(\edb_top_inst/n3639 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5171 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__5172  (.I0(\edb_top_inst/n3636 ), .I1(\edb_top_inst/n3635 ), 
            .I2(\edb_top_inst/n3637 ), .I3(\edb_top_inst/n3639 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5172 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__5173  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/n3630 ), 
            .I2(\edb_top_inst/n3596 ), .I3(\edb_top_inst/n3597 ), .O(\edb_top_inst/n3640 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5173 .LUTMASK = 16'hbe00;
    EFX_LUT4 \edb_top_inst/LUT__5174  (.I0(\edb_top_inst/n3584 ), .I1(\edb_top_inst/n3564 ), 
            .I2(\edb_top_inst/n3591 ), .O(\edb_top_inst/n3641 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5174 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__5175  (.I0(\edb_top_inst/n3538 ), .I1(\edb_top_inst/n3558 ), 
            .I2(\edb_top_inst/n3641 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3642 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5175 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__5176  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3643 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5176 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__5177  (.I0(\edb_top_inst/n3599 ), .I1(\edb_top_inst/n3591 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3644 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5177 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__5178  (.I0(\edb_top_inst/n3620 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3644 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n3645 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5178 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__5179  (.I0(\edb_top_inst/n3620 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3626 ), .O(\edb_top_inst/n3646 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5179 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__5180  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n3624 ), .I2(\edb_top_inst/n3645 ), .I3(\edb_top_inst/n3646 ), 
            .O(\edb_top_inst/n3647 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5180 .LUTMASK = 16'h00fe;
    EFX_LUT4 \edb_top_inst/LUT__5181  (.I0(\edb_top_inst/n3642 ), .I1(\edb_top_inst/n3640 ), 
            .I2(\edb_top_inst/n3643 ), .I3(\edb_top_inst/n3647 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5181 .LUTMASK = 16'h10ff;
    EFX_LUT4 \edb_top_inst/LUT__5182  (.I0(\edb_top_inst/la0/la_biu_inst/n374 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
            .O(\edb_top_inst/ceg_net348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5182 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__5183  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5183 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5184  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I2(\edb_top_inst/n3259 ), 
            .O(\edb_top_inst/n3648 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5184 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5185  (.I0(\edb_top_inst/n3594 ), .I1(\edb_top_inst/n3648 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n2043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5185 .LUTMASK = 16'h7777;
    EFX_LUT4 \edb_top_inst/LUT__5186  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5186 .LUTMASK = 16'h05fc;
    EFX_LUT4 \edb_top_inst/LUT__5187  (.I0(\edb_top_inst/la0/la_biu_inst/n2043 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n3649 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5187 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5188  (.I0(\edb_top_inst/n3517 ), .I1(\edb_top_inst/n3649 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5188 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5189  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I2(\edb_top_inst/n3259 ), 
            .I3(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5189 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__5190  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5190 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__5191  (.I0(\edb_top_inst/n3649 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/ceg_net355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5191 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5192  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .I1(\edb_top_inst/n3260 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5192 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__5193  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[15] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5193 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5194  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[16] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5194 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5195  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[17] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5195 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5196  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[18] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5196 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5197  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[19] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5197 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5198  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[20] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5198 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5199  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[21] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5199 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5200  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[22] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5200 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5201  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[23] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5201 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5202  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[24] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5202 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5203  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[25] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5203 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5204  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[26] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5204 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5205  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[12] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[27] ), .I2(\edb_top_inst/n3260 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5205 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5206  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I1(\edb_top_inst/n3511 ), .O(\edb_top_inst/n3650 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5206 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5207  (.I0(\edb_top_inst/n3495 ), .I1(\edb_top_inst/n3650 ), 
            .O(\edb_top_inst/n3651 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5207 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5208  (.I0(\edb_top_inst/n3549 ), .I1(\edb_top_inst/n3550 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .I3(\edb_top_inst/n3651 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5208 .LUTMASK = 16'hffe0;
    EFX_LUT4 \edb_top_inst/LUT__5209  (.I0(\edb_top_inst/n3493 ), .I1(\edb_top_inst/n3490 ), 
            .O(\edb_top_inst/n3652 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5209 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5210  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3653 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5210 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__5211  (.I0(\edb_top_inst/n3653 ), .I1(\edb_top_inst/n3499 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I3(\edb_top_inst/n3652 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5211 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__5212  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/n3498 ), 
            .I3(\edb_top_inst/n3490 ), .O(\edb_top_inst/n3654 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5212 .LUTMASK = 16'hfe00;
    EFX_LUT4 \edb_top_inst/LUT__5213  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3655 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5213 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5214  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/n3655 ), 
            .I3(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3656 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5214 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__5215  (.I0(\edb_top_inst/n3656 ), .I1(\edb_top_inst/n3499 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I3(\edb_top_inst/n3654 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5215 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__5216  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/n3490 ), 
            .O(\edb_top_inst/n3657 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5216 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__5217  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3658 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5217 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5218  (.I0(\edb_top_inst/n3658 ), .I1(\edb_top_inst/n3655 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3659 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5218 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5219  (.I0(\edb_top_inst/n3659 ), .I1(\edb_top_inst/n3499 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I3(\edb_top_inst/n3657 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5219 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__5220  (.I0(\edb_top_inst/n3504 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[3] ), .I3(\edb_top_inst/n3490 ), 
            .O(\edb_top_inst/n3660 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5220 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__5221  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5221 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5222  (.I0(\edb_top_inst/n3661 ), .I1(\edb_top_inst/n3658 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3662 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5222 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5223  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I1(\edb_top_inst/n3504 ), .I2(\edb_top_inst/n3662 ), .I3(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3663 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5223 .LUTMASK = 16'h77f0;
    EFX_LUT4 \edb_top_inst/LUT__5224  (.I0(\edb_top_inst/n3663 ), .I1(\edb_top_inst/n3495 ), 
            .O(\edb_top_inst/n3664 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5224 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5225  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(\edb_top_inst/n3660 ), .I2(\edb_top_inst/n3664 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5225 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5226  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3665 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5226 .LUTMASK = 16'h0708;
    EFX_LUT4 \edb_top_inst/LUT__5227  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5227 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5228  (.I0(\edb_top_inst/n3666 ), .I1(\edb_top_inst/n3661 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3667 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5228 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5229  (.I0(\edb_top_inst/n3667 ), .I1(\edb_top_inst/n3653 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3495 ), 
            .O(\edb_top_inst/n3668 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5229 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__5230  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(\edb_top_inst/n3665 ), .I2(\edb_top_inst/n3668 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5230 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5231  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3669 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5231 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__5232  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3670 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5232 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5233  (.I0(\edb_top_inst/n3670 ), .I1(\edb_top_inst/n3666 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3671 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5233 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5234  (.I0(\edb_top_inst/n3671 ), .I1(\edb_top_inst/n3656 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3495 ), 
            .O(\edb_top_inst/n3672 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5234 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__5235  (.I0(\edb_top_inst/n3669 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I2(\edb_top_inst/n3665 ), .I3(\edb_top_inst/n3672 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5235 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5236  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/n3665 ), 
            .O(\edb_top_inst/n3673 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5236 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__5237  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3674 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5237 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5238  (.I0(\edb_top_inst/n3674 ), .I1(\edb_top_inst/n3670 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3675 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5238 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5239  (.I0(\edb_top_inst/n3675 ), .I1(\edb_top_inst/n3659 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3495 ), 
            .O(\edb_top_inst/n3676 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5239 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__5240  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I1(\edb_top_inst/n3673 ), .I2(\edb_top_inst/n3676 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5240 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5241  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5241 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5242  (.I0(\edb_top_inst/n3677 ), .I1(\edb_top_inst/n3674 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3678 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5242 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5243  (.I0(\edb_top_inst/n3678 ), .I1(\edb_top_inst/n3662 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3679 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5243 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5244  (.I0(\edb_top_inst/n3679 ), .I1(\edb_top_inst/n3650 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3680 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5244 .LUTMASK = 16'h0c05;
    EFX_LUT4 \edb_top_inst/LUT__5245  (.I0(\edb_top_inst/n3511 ), .I1(\edb_top_inst/n3673 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I3(\edb_top_inst/n3680 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5245 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5246  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3681 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5246 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__5247  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5247 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5248  (.I0(\edb_top_inst/n3682 ), .I1(\edb_top_inst/n3677 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5248 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5249  (.I0(\edb_top_inst/n3683 ), .I1(\edb_top_inst/n3653 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5249 .LUTMASK = 16'h0c05;
    EFX_LUT4 \edb_top_inst/LUT__5250  (.I0(\edb_top_inst/n3667 ), .I1(\edb_top_inst/n3681 ), 
            .I2(\edb_top_inst/n3684 ), .I3(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5250 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__5251  (.I0(\edb_top_inst/n3496 ), .I1(\edb_top_inst/n3673 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I3(\edb_top_inst/n3685 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5251 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5252  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5252 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__5253  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5253 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5254  (.I0(\edb_top_inst/n3687 ), .I1(\edb_top_inst/n3682 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5254 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5255  (.I0(\edb_top_inst/n3688 ), .I1(\edb_top_inst/n3656 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5255 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__5256  (.I0(\edb_top_inst/n3671 ), .I1(\edb_top_inst/n3681 ), 
            .I2(\edb_top_inst/n3689 ), .I3(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5256 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__5257  (.I0(\edb_top_inst/n3686 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I2(\edb_top_inst/n3665 ), .I3(\edb_top_inst/n3690 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5257 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5258  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5258 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5259  (.I0(\edb_top_inst/n3691 ), .I1(\edb_top_inst/n3687 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5259 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5260  (.I0(\edb_top_inst/n3692 ), .I1(\edb_top_inst/n3659 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5260 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__5261  (.I0(\edb_top_inst/n3675 ), .I1(\edb_top_inst/n3681 ), 
            .I2(\edb_top_inst/n3693 ), .I3(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5261 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__5262  (.I0(\edb_top_inst/n3548 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] ), 
            .I2(\edb_top_inst/n3694 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5262 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5263  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5263 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__5264  (.I0(\edb_top_inst/n3695 ), .I1(\edb_top_inst/n3691 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5264 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5265  (.I0(\edb_top_inst/n3696 ), .I1(\edb_top_inst/n3678 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5265 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__5266  (.I0(\edb_top_inst/n3697 ), .I1(\edb_top_inst/n3663 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5266 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__5267  (.I0(\edb_top_inst/n3549 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12] ), 
            .I2(\edb_top_inst/n3698 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5267 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5268  (.I0(\edb_top_inst/n3549 ), .I1(\edb_top_inst/n3550 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .I3(\edb_top_inst/n3651 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5268 .LUTMASK = 16'hffe0;
    EFX_LUT4 \edb_top_inst/LUT__5269  (.I0(\edb_top_inst/n3653 ), .I1(\edb_top_inst/n3499 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I3(\edb_top_inst/n3652 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5269 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__5270  (.I0(\edb_top_inst/n3656 ), .I1(\edb_top_inst/n3499 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I3(\edb_top_inst/n3654 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5270 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__5271  (.I0(\edb_top_inst/n3659 ), .I1(\edb_top_inst/n3499 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I3(\edb_top_inst/n3657 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5271 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__5272  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(\edb_top_inst/n3660 ), .I2(\edb_top_inst/n3664 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5272 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5273  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(\edb_top_inst/n3665 ), .I2(\edb_top_inst/n3668 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5273 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5274  (.I0(\edb_top_inst/n3669 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I2(\edb_top_inst/n3665 ), .I3(\edb_top_inst/n3672 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5274 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5275  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I1(\edb_top_inst/n3673 ), .I2(\edb_top_inst/n3676 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5275 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5276  (.I0(\edb_top_inst/n3511 ), .I1(\edb_top_inst/n3673 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I3(\edb_top_inst/n3680 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5276 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5277  (.I0(\edb_top_inst/n3496 ), .I1(\edb_top_inst/n3673 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I3(\edb_top_inst/n3685 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5277 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5278  (.I0(\edb_top_inst/n3686 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I2(\edb_top_inst/n3665 ), .I3(\edb_top_inst/n3690 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5278 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__5279  (.I0(\edb_top_inst/n3548 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] ), 
            .I2(\edb_top_inst/n3694 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5279 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5280  (.I0(\edb_top_inst/n3549 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12] ), 
            .I2(\edb_top_inst/n3698 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5280 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__5281  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .I2(\edb_top_inst/la0/module_state[0] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3699 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcc53, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5281 .LUTMASK = 16'hcc53;
    EFX_LUT4 \edb_top_inst/LUT__5282  (.I0(\edb_top_inst/n3699 ), .I1(jtag_inst2_UPDATE), 
            .I2(\edb_top_inst/edb_user_dr[81] ), .I3(jtag_inst2_SEL), .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5282 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__5283  (.I0(jtag_inst2_SEL), .I1(jtag_inst2_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5283 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__5284  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[1] ), .O(\edb_top_inst/n3096 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5284 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__5289  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5289 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5293  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5293 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5294  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i2_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5294 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5295  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5295 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5296  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5296 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5297  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5297 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5298  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5298 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5299  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5299 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5300  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5300 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5301  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5301 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5302  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5302 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5303  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i24_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5303 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5304  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5304 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5305  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5305 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5306  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5306 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5307  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5307 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5308  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5308 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5309  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i3_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5309 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5310  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5310 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5311  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5311 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5312  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i6_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5312 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5313  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i7_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5313 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5314  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5314 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5315  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5315 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5316  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5316 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5317  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5317 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5318  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5318 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5319  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5319 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5320  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5320 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5321  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5321 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5322  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5322 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5323  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5323 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5324  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i1_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5324 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__5325  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__5325 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4316  (.I0(\edb_top_inst/la0/crc_data_out[16] ), 
            .I1(\edb_top_inst/edb_user_dr[66] ), .I2(\edb_top_inst/la0/crc_data_out[23] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n3115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4316 .LUTMASK = 16'h9009;
    EFX_RAM10 \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram  (.WCLK(1'b0), 
            .RCLK(iBCLK), .WCLKE(1'b0), .RE(1'b1), .RST(1'b0), .WADDREN(1'b0), 
            .RADDREN(1'b1), .WE({2'b00}), .WADDR({10'b0000000000}), .RADDR({\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[1] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[0] }), .RDATA({\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=8, WRITE_WIDTH=8, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="NONE", INIT_0=256'h1F24AD230422DC211D201B1F1C1E001D001CAD1B041A3419E71838160115C0D6, INIT_1=256'hC0962856005508481041772F1B2E7C2D082CAD2B042A00290028352701262425, INIT_2=256'h007F00F980FEE0FDE09A01DFD0E0C0D660BA06AFA4A3A4A2619D309CE09A0398, INIT_3=256'h0000000000000000000000000000000000000000000000000000104101E20094, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .READ_WIDTH = 8;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WRITE_WIDTH = 8;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RESET_OUTREG = "NONE";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_0 = 256'h1F24AD230422DC211D201B1F1C1E001D001CAD1B041A3419E71838160115C0D6;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1 = 256'hC0962856005508481041772F1B2E7C2D082CAD2B042A00290028352701262425;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_2 = 256'h007F00F980FEE0FDE09A01DFD0E0C0D660BA06AFA4A3A4A2619D309CE09A0398;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000104101E20094;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .OUTPUT_REG = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_ADD \edb_top_inst/la0/add_91/i1  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/n1224 ), .CI(1'b0), .O(\edb_top_inst/n59 ), 
            .CO(\edb_top_inst/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i2  (.I0(\edb_top_inst/la0/bit_count[1] ), 
            .I1(\edb_top_inst/la0/bit_count[0] ), .CI(1'b0), .O(\edb_top_inst/n61 ), 
            .CO(\edb_top_inst/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_100/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n662 ), .CO(\edb_top_inst/n663 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n664 ), .CO(\edb_top_inst/n665 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .CI(1'b0), 
            .CO(\edb_top_inst/n666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[0] ), .CI(1'b0), .CO(\edb_top_inst/n667 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(1'b1), .CI(n10448), .O(\edb_top_inst/n877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4701)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(1'b1), .CI(n10449), .O(\edb_top_inst/n878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4687)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i14  (.I0(\edb_top_inst/la0/la_sample_cnt[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/n881 ), .O(\edb_top_inst/n879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13  (.I0(\edb_top_inst/la0/la_sample_cnt[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n883 ), .O(\edb_top_inst/n880 ), 
            .CO(\edb_top_inst/n881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n885 ), .O(\edb_top_inst/n882 ), 
            .CO(\edb_top_inst/n883 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n887 ), .O(\edb_top_inst/n884 ), 
            .CO(\edb_top_inst/n885 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n889 ), .O(\edb_top_inst/n886 ), 
            .CO(\edb_top_inst/n887 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n891 ), .O(\edb_top_inst/n888 ), 
            .CO(\edb_top_inst/n889 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n893 ), .O(\edb_top_inst/n890 ), 
            .CO(\edb_top_inst/n891 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n895 ), .O(\edb_top_inst/n892 ), 
            .CO(\edb_top_inst/n893 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n897 ), .O(\edb_top_inst/n894 ), 
            .CO(\edb_top_inst/n895 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n899 ), .O(\edb_top_inst/n896 ), 
            .CO(\edb_top_inst/n897 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n901 ), .O(\edb_top_inst/n898 ), 
            .CO(\edb_top_inst/n899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n667 ), .O(\edb_top_inst/n900 ), 
            .CO(\edb_top_inst/n901 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4703)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i14  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/n904 ), .O(\edb_top_inst/n902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n906 ), .O(\edb_top_inst/n903 ), 
            .CO(\edb_top_inst/n904 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n908 ), .O(\edb_top_inst/n905 ), 
            .CO(\edb_top_inst/n906 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n910 ), .O(\edb_top_inst/n907 ), 
            .CO(\edb_top_inst/n908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n912 ), .O(\edb_top_inst/n909 ), 
            .CO(\edb_top_inst/n910 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n914 ), .O(\edb_top_inst/n911 ), 
            .CO(\edb_top_inst/n912 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n916 ), .O(\edb_top_inst/n913 ), 
            .CO(\edb_top_inst/n914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n918 ), .O(\edb_top_inst/n915 ), 
            .CO(\edb_top_inst/n916 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n920 ), .O(\edb_top_inst/n917 ), 
            .CO(\edb_top_inst/n918 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n922 ), .O(\edb_top_inst/n919 ), 
            .CO(\edb_top_inst/n920 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n924 ), .O(\edb_top_inst/n921 ), 
            .CO(\edb_top_inst/n922 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n666 ), .O(\edb_top_inst/n923 ), 
            .CO(\edb_top_inst/n924 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4689)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i13  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n954 ), .O(\edb_top_inst/n951 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n956 ), .O(\edb_top_inst/n953 ), 
            .CO(\edb_top_inst/n954 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n958 ), .O(\edb_top_inst/n955 ), 
            .CO(\edb_top_inst/n956 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n960 ), .O(\edb_top_inst/n957 ), 
            .CO(\edb_top_inst/n958 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n962 ), .O(\edb_top_inst/n959 ), 
            .CO(\edb_top_inst/n960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n964 ), .O(\edb_top_inst/n961 ), 
            .CO(\edb_top_inst/n962 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n966 ), .O(\edb_top_inst/n963 ), 
            .CO(\edb_top_inst/n964 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n968 ), .O(\edb_top_inst/n965 ), 
            .CO(\edb_top_inst/n966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n970 ), .O(\edb_top_inst/n967 ), 
            .CO(\edb_top_inst/n968 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n972 ), .O(\edb_top_inst/n969 ), 
            .CO(\edb_top_inst/n970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n665 ), .O(\edb_top_inst/n971 ), 
            .CO(\edb_top_inst/n972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4682)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i13  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n977 ), .O(\edb_top_inst/n974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n979 ), .O(\edb_top_inst/n976 ), 
            .CO(\edb_top_inst/n977 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n982 ), .O(\edb_top_inst/n978 ), 
            .CO(\edb_top_inst/n979 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n985 ), .O(\edb_top_inst/n981 ), 
            .CO(\edb_top_inst/n982 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n987 ), .O(\edb_top_inst/n984 ), 
            .CO(\edb_top_inst/n985 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n989 ), .O(\edb_top_inst/n986 ), 
            .CO(\edb_top_inst/n987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n991 ), .O(\edb_top_inst/n988 ), 
            .CO(\edb_top_inst/n989 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n993 ), .O(\edb_top_inst/n990 ), 
            .CO(\edb_top_inst/n991 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n995 ), .O(\edb_top_inst/n992 ), 
            .CO(\edb_top_inst/n993 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n997 ), .O(\edb_top_inst/n994 ), 
            .CO(\edb_top_inst/n995 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n663 ), .O(\edb_top_inst/n996 ), 
            .CO(\edb_top_inst/n997 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4678)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i13  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1000 ), .O(\edb_top_inst/n998 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1002 ), .O(\edb_top_inst/n999 ), 
            .CO(\edb_top_inst/n1000 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1004 ), .O(\edb_top_inst/n1001 ), 
            .CO(\edb_top_inst/n1002 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1006 ), .O(\edb_top_inst/n1003 ), 
            .CO(\edb_top_inst/n1004 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1008 ), .O(\edb_top_inst/n1005 ), 
            .CO(\edb_top_inst/n1006 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1010 ), .O(\edb_top_inst/n1007 ), 
            .CO(\edb_top_inst/n1008 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1012 ), .O(\edb_top_inst/n1009 ), 
            .CO(\edb_top_inst/n1010 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1014 ), .O(\edb_top_inst/n1011 ), 
            .CO(\edb_top_inst/n1012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1016 ), .O(\edb_top_inst/n1013 ), 
            .CO(\edb_top_inst/n1014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1018 ), .O(\edb_top_inst/n1015 ), 
            .CO(\edb_top_inst/n1016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1020 ), .O(\edb_top_inst/n1017 ), 
            .CO(\edb_top_inst/n1018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .CI(1'b0), 
            .O(\edb_top_inst/n1019 ), .CO(\edb_top_inst/n1020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4671)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i6  (.I0(\edb_top_inst/la0/bit_count[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1023 ), .O(\edb_top_inst/n1021 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_100/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i5  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1025 ), .O(\edb_top_inst/n1022 ), 
            .CO(\edb_top_inst/n1023 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_100/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i4  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1027 ), .O(\edb_top_inst/n1024 ), 
            .CO(\edb_top_inst/n1025 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_100/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i3  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n62 ), .O(\edb_top_inst/n1026 ), 
            .CO(\edb_top_inst/n1027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3749)
    defparam \edb_top_inst/la0/add_100/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i28  (.I0(\edb_top_inst/la0/address_counter[27] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1038 ), .O(\edb_top_inst/n1035 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i28 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i27  (.I0(\edb_top_inst/la0/address_counter[26] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1040 ), .O(\edb_top_inst/n1037 ), 
            .CO(\edb_top_inst/n1038 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i27 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i26  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1042 ), .O(\edb_top_inst/n1039 ), 
            .CO(\edb_top_inst/n1040 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i26 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i25  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1044 ), .O(\edb_top_inst/n1041 ), 
            .CO(\edb_top_inst/n1042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i24  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1046 ), .O(\edb_top_inst/n1043 ), 
            .CO(\edb_top_inst/n1044 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i23  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1048 ), .O(\edb_top_inst/n1045 ), 
            .CO(\edb_top_inst/n1046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i22  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1050 ), .O(\edb_top_inst/n1047 ), 
            .CO(\edb_top_inst/n1048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i21  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1052 ), .O(\edb_top_inst/n1049 ), 
            .CO(\edb_top_inst/n1050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i20  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1054 ), .O(\edb_top_inst/n1051 ), 
            .CO(\edb_top_inst/n1052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i19  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1056 ), .O(\edb_top_inst/n1053 ), 
            .CO(\edb_top_inst/n1054 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i18  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1058 ), .O(\edb_top_inst/n1055 ), 
            .CO(\edb_top_inst/n1056 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i17  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1060 ), .O(\edb_top_inst/n1057 ), 
            .CO(\edb_top_inst/n1058 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i16  (.I0(\edb_top_inst/la0/address_counter[15] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1062 ), .O(\edb_top_inst/n1059 ), 
            .CO(\edb_top_inst/n1060 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i15  (.I0(\edb_top_inst/la0/address_counter[14] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1064 ), .O(\edb_top_inst/n1061 ), 
            .CO(\edb_top_inst/n1062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i14  (.I0(\edb_top_inst/la0/address_counter[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1066 ), .O(\edb_top_inst/n1063 ), 
            .CO(\edb_top_inst/n1064 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i13  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1068 ), .O(\edb_top_inst/n1065 ), 
            .CO(\edb_top_inst/n1066 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i12  (.I0(\edb_top_inst/la0/address_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1070 ), .O(\edb_top_inst/n1067 ), 
            .CO(\edb_top_inst/n1068 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i11  (.I0(\edb_top_inst/la0/address_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1072 ), .O(\edb_top_inst/n1069 ), 
            .CO(\edb_top_inst/n1070 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i10  (.I0(\edb_top_inst/la0/address_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1074 ), .O(\edb_top_inst/n1071 ), 
            .CO(\edb_top_inst/n1072 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i9  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1076 ), .O(\edb_top_inst/n1073 ), 
            .CO(\edb_top_inst/n1074 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i8  (.I0(\edb_top_inst/la0/address_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1078 ), .O(\edb_top_inst/n1075 ), 
            .CO(\edb_top_inst/n1076 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i7  (.I0(\edb_top_inst/la0/address_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1080 ), .O(\edb_top_inst/n1077 ), 
            .CO(\edb_top_inst/n1078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i6  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1082 ), .O(\edb_top_inst/n1079 ), 
            .CO(\edb_top_inst/n1080 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i5  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1084 ), .O(\edb_top_inst/n1081 ), 
            .CO(\edb_top_inst/n1082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i4  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/n3090 ), .CI(\edb_top_inst/n1086 ), .O(\edb_top_inst/n1083 ), 
            .CO(\edb_top_inst/n1084 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i3  (.I0(\edb_top_inst/la0/address_counter[2] ), 
            .I1(\edb_top_inst/n3093 ), .CI(\edb_top_inst/n1088 ), .O(\edb_top_inst/n1085 ), 
            .CO(\edb_top_inst/n1086 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i2  (.I0(\edb_top_inst/la0/address_counter[1] ), 
            .I1(\edb_top_inst/n3096 ), .CI(\edb_top_inst/n60 ), .O(\edb_top_inst/n1087 ), 
            .CO(\edb_top_inst/n1088 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3722)
    defparam \edb_top_inst/la0/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i13  (.I0(\edb_top_inst/la0/address_counter[27] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1099 ), .O(\edb_top_inst/n1096 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i12  (.I0(\edb_top_inst/la0/address_counter[26] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1101 ), .O(\edb_top_inst/n1098 ), 
            .CO(\edb_top_inst/n1099 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i11  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1103 ), .O(\edb_top_inst/n1100 ), 
            .CO(\edb_top_inst/n1101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i10  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1105 ), .O(\edb_top_inst/n1102 ), 
            .CO(\edb_top_inst/n1103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i9  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1107 ), .O(\edb_top_inst/n1104 ), 
            .CO(\edb_top_inst/n1105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i8  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1109 ), .O(\edb_top_inst/n1106 ), 
            .CO(\edb_top_inst/n1107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i7  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1111 ), .O(\edb_top_inst/n1108 ), 
            .CO(\edb_top_inst/n1109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i6  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1116 ), .O(\edb_top_inst/n1110 ), 
            .CO(\edb_top_inst/n1111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i5  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1118 ), .O(\edb_top_inst/n1115 ), 
            .CO(\edb_top_inst/n1116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i4  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1120 ), .O(\edb_top_inst/n1117 ), 
            .CO(\edb_top_inst/n1118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i3  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1203 ), .O(\edb_top_inst/n1119 ), 
            .CO(\edb_top_inst/n1120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i2  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(\edb_top_inst/la0/address_counter[15] ), .CI(1'b0), .O(\edb_top_inst/n1202 ), 
            .CO(\edb_top_inst/n1203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/kimura/workspace/ProjectFolder/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_90/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i2 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__13847 (.I0(n10054), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .O(\MCsiRxController/MCsi2Decoder/select_39/Select_0/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13847.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13848 (.I0(oTestPort[25]), .I1(MipiDphyRx1_RX_SYNC_HS_LAN1), 
            .O(\MCsiRxController/MCsi2Decoder/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__13848.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__13849 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .O(n10055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13849.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13850 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[10] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10] ), 
            .O(n10056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13850.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13851 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .O(n10057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13851.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13852 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .O(n10058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13852.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13853 (.I0(n10055), .I1(n10056), .I2(n10057), .I3(n10058), 
            .O(n10059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13853.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13854 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .O(n10060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13854.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13855 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I2(n10059), .I3(n10060), .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6fff */ ;
    defparam LUT__13855.LUTMASK = 16'h6fff;
    EFX_LUT4 LUT__13856 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .O(n10061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13856.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13857 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(n10062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13857.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13858 (.I0(n10061), .I1(n10062), .O(n10063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13858.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13859 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .O(n10064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__13859.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__13860 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[10] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] ), 
            .O(n10065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13860.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13861 (.I0(n10065), .I1(n10063), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .O(n10066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd73d */ ;
    defparam LUT__13861.LUTMASK = 16'hd73d;
    EFX_LUT4 LUT__13862 (.I0(n10064), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I2(n10063), .I3(n10066), .O(n10067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__13862.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__13863 (.I0(n10061), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(n10068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13863.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13864 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(n10069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13864.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13865 (.I0(n10069), .I1(n10061), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(n10070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__13865.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__13866 (.I0(n10070), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .I3(n10068), .O(n10071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1441 */ ;
    defparam LUT__13866.LUTMASK = 16'h1441;
    EFX_LUT4 LUT__13867 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .O(n10072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13867.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13868 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n10073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__13868.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__13869 (.I0(n10073), .I1(n10072), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .O(n10074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha333 */ ;
    defparam LUT__13869.LUTMASK = 16'ha333;
    EFX_LUT4 LUT__13870 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .O(n10075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13870.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13871 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .O(n10076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13871.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13872 (.I0(n10076), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I3(n10075), .O(n10077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800 */ ;
    defparam LUT__13872.LUTMASK = 16'h1800;
    EFX_LUT4 LUT__13873 (.I0(n10074), .I1(n10071), .I2(n10077), .O(n10078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13873.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13874 (.I0(n10061), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .O(n10079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13874.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13875 (.I0(n10079), .I1(n10062), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .O(n10080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13875.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13876 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n10081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13876.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13877 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(n10082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13877.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13878 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(n10081), .I2(n10082), .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .O(n10083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__13878.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__13879 (.I0(n10069), .I1(n10079), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(n10084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__13879.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__13880 (.I0(n10080), .I1(n10064), .I2(n10083), .I3(n10084), 
            .O(n10085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__13880.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__13881 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(n10086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__13881.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__13882 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .O(n10087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13882.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13883 (.I0(n10086), .I1(n10087), .I2(n10068), .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .O(n10088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccc */ ;
    defparam LUT__13883.LUTMASK = 16'h5ccc;
    EFX_LUT4 LUT__13884 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .O(n10089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__13884.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__13885 (.I0(n10082), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n10090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13885.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13886 (.I0(n10089), .I1(n10090), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .O(n10091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1441 */ ;
    defparam LUT__13886.LUTMASK = 16'h1441;
    EFX_LUT4 LUT__13887 (.I0(n10080), .I1(n10065), .I2(n10088), .I3(n10091), 
            .O(n10092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__13887.LUTMASK = 16'he000;
    EFX_LUT4 LUT__13888 (.I0(n10085), .I1(n10092), .I2(n10067), .I3(n10078), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qFullAllmost )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__13888.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__13889 (.I0(n10069), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I3(n10065), .O(n10093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100 */ ;
    defparam LUT__13889.LUTMASK = 16'h4100;
    EFX_LUT4 LUT__13890 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I2(n10076), .I3(n10075), .O(n10094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__13890.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__13891 (.I0(n10093), .I1(n10094), .I2(n10087), .I3(n10072), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__13891.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__13892 (.I0(\MCsiRxController/MCsi2Decoder/wFtiEmp[0] ), 
            .I1(wCdcFifoFull), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n21 ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13892.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13893 (.I0(\wHsDatatype[2] ), .I1(\wHsDatatype[3] ), .I2(\wHsDatatype[4] ), 
            .I3(\wHsDatatype[5] ), .O(n10095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__13893.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__13894 (.I0(n10095), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I3(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .O(n10096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff3 */ ;
    defparam LUT__13894.LUTMASK = 16'heff3;
    EFX_LUT4 LUT__13895 (.I0(n10096), .I1(rSRST), .I2(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .O(\MCsiRxController/MCsi2Decoder/n640 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__13895.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__13896 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .I3(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .O(\MCsiRxController/MCsi2Decoder/n659 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800 */ ;
    defparam LUT__13896.LUTMASK = 16'h1800;
    EFX_LUT4 LUT__13897 (.I0(\wHsWordCnt[12] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .O(n10097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13897.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13898 (.I0(\wHsWordCnt[14] ), .I1(n10097), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] ), 
            .I3(\wHsWordCnt[13] ), .O(n10098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7e */ ;
    defparam LUT__13898.LUTMASK = 16'heb7e;
    EFX_LUT4 LUT__13899 (.I0(\wHsWordCnt[1] ), .I1(\wHsWordCnt[2] ), .I2(\wHsWordCnt[3] ), 
            .I3(\wHsWordCnt[4] ), .O(n10099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13899.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13900 (.I0(\wHsWordCnt[5] ), .I1(\wHsWordCnt[6] ), .I2(\wHsWordCnt[7] ), 
            .I3(\wHsWordCnt[8] ), .O(n10100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13900.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13901 (.I0(\wHsWordCnt[9] ), .I1(\wHsWordCnt[10] ), .I2(n10099), 
            .I3(n10100), .O(n10101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13901.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13902 (.I0(\wHsWordCnt[14] ), .I1(\wHsWordCnt[13] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] ), 
            .I3(\wHsWordCnt[11] ), .O(n10102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100 */ ;
    defparam LUT__13902.LUTMASK = 16'h4100;
    EFX_LUT4 LUT__13903 (.I0(n10098), .I1(n10101), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I3(n10102), .O(n10103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00be */ ;
    defparam LUT__13903.LUTMASK = 16'h00be;
    EFX_LUT4 LUT__13904 (.I0(\wHsWordCnt[12] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), .O(n10104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__13904.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__13905 (.I0(n10099), .I1(n10100), .O(n10105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13905.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13906 (.I0(\wHsWordCnt[9] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] ), 
            .O(n10106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13906.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13907 (.I0(n10101), .I1(n10104), .I2(n10105), .I3(n10106), 
            .O(n10107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7007 */ ;
    defparam LUT__13907.LUTMASK = 16'h7007;
    EFX_LUT4 LUT__13908 (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), 
            .I1(\wHsWordCnt[2] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] ), 
            .I3(\wHsWordCnt[1] ), .O(n10108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7 */ ;
    defparam LUT__13908.LUTMASK = 16'hbed7;
    EFX_LUT4 LUT__13909 (.I0(\wHsWordCnt[11] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I2(\wHsWordCnt[12] ), .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .O(n10109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bb0 */ ;
    defparam LUT__13909.LUTMASK = 16'h0bb0;
    EFX_LUT4 LUT__13910 (.I0(n10108), .I1(n10109), .I2(\wHsWordCnt[15] ), 
            .I3(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), .O(n10110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13910.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13911 (.I0(n10103), .I1(n10107), .I2(n10110), .O(n10111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13911.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13912 (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I1(\wHsWordCnt[11] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] ), 
            .I3(\wHsWordCnt[10] ), .O(n10112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40f */ ;
    defparam LUT__13912.LUTMASK = 16'hf40f;
    EFX_LUT4 LUT__13913 (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I1(\wHsWordCnt[11] ), .I2(\wHsWordCnt[10] ), .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] ), 
            .O(n10113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b */ ;
    defparam LUT__13913.LUTMASK = 16'hb00b;
    EFX_LUT4 LUT__13914 (.I0(n10112), .I1(n10113), .I2(\wHsWordCnt[9] ), 
            .I3(n10105), .O(n10114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5cc */ ;
    defparam LUT__13914.LUTMASK = 16'hc5cc;
    EFX_LUT4 LUT__13915 (.I0(\wHsWordCnt[5] ), .I1(\wHsWordCnt[6] ), .I2(n10099), 
            .O(n10115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13915.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13916 (.I0(\wHsWordCnt[8] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] ), 
            .O(n10116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13916.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13917 (.I0(n10116), .I1(n10115), .I2(\wHsWordCnt[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] ), .O(n10117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__13917.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__13918 (.I0(\wHsWordCnt[1] ), .I1(\wHsWordCnt[2] ), .O(n10118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13918.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13919 (.I0(\wHsWordCnt[4] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] ), 
            .O(n10119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13919.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13920 (.I0(n10119), .I1(n10118), .I2(\wHsWordCnt[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] ), .O(n10120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__13920.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__13921 (.I0(\wHsWordCnt[6] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] ), 
            .O(n10121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13921.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13922 (.I0(n10121), .I1(n10099), .I2(\wHsWordCnt[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] ), .O(n10122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__13922.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__13923 (.I0(n10117), .I1(n10120), .I2(n10122), .I3(n10114), 
            .O(n10123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13923.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13924 (.I0(n10123), .I1(n10111), .I2(rSRST), .O(\MCsiRxController/MCsi2Decoder/qLineCntRst )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__13924.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__13925 (.I0(n10095), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .I3(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .O(n10124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb0f */ ;
    defparam LUT__13925.LUTMASK = 16'hfb0f;
    EFX_LUT4 LUT__13927 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .I1(n10123), 
            .I2(n10111), .I3(n10124), .O(\MCsiRxController/MCsi2Decoder/select_39/Select_2/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__13927.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__13845 (.I0(pll_inst1_LOCKED), .I1(pll_inst2_LOCKED), .O(oLed[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13845.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13928 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .O(\MCsiRxController/MCsi2Decoder/equal_30/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__13928.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__13929 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), .O(\MCsiRxController/MCsi2Decoder/equal_31/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__13929.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__13930 (.I0(\MCsiRxController/MCsi2Decoder/equal_30/n8 ), 
            .I1(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), .I2(\MCsiRxController/MCsi2Decoder/equal_31/n8 ), 
            .O(\MCsiRxController/MCsi2Decoder/select_39/Select_1/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__13930.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__13931 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13931.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13932 (.I0(n10082), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13932.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13933 (.I0(n10082), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13933.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13934 (.I0(n10090), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13934.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13935 (.I0(n10079), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13935.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13936 (.I0(n10079), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13936.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13937 (.I0(n10068), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13937.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13938 (.I0(n10063), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13938.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13939 (.I0(n10080), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n305 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13939.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13940 (.I0(n10080), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[10] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13940.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13941 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .O(n10126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__13941.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__13942 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), .O(n10127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13942.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13943 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] ), .O(n10128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13943.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13944 (.I0(n10128), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), .O(n10129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__13944.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__13945 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), .O(n10130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13945.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13946 (.I0(n10127), .I1(n10126), .I2(n10129), .I3(n10130), 
            .O(n10131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13946.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13947 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), .O(n10132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13947.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13948 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), .I2(n10131), 
            .I3(n10132), .O(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6fff */ ;
    defparam LUT__13948.LUTMASK = 16'h6fff;
    EFX_LUT4 LUT__13949 (.I0(\MCsiRxController/wFtiEmp[0] ), .I1(wVideofull), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__13949.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__13950 (.I0(n10126), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .I3(n10127), 
            .O(n10133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef54 */ ;
    defparam LUT__13950.LUTMASK = 16'hef54;
    EFX_LUT4 LUT__13951 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), .I2(n10126), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), .O(n10134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e9f */ ;
    defparam LUT__13951.LUTMASK = 16'h7e9f;
    EFX_LUT4 LUT__13952 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .O(n10135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13952.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13953 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I1(n10128), .I2(n10135), .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .O(n10136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde */ ;
    defparam LUT__13953.LUTMASK = 16'hbdde;
    EFX_LUT4 LUT__13954 (.I0(n10136), .I1(n10129), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(n10137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa3f */ ;
    defparam LUT__13954.LUTMASK = 16'hfa3f;
    EFX_LUT4 LUT__13955 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), 
            .I3(n10127), .O(n10138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef51 */ ;
    defparam LUT__13955.LUTMASK = 16'hef51;
    EFX_LUT4 LUT__13956 (.I0(n10126), .I1(n10138), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), .O(n10139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0230 */ ;
    defparam LUT__13956.LUTMASK = 16'h0230;
    EFX_LUT4 LUT__13957 (.I0(n10136), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(n10140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__13957.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__13958 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), .O(n10141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__13958.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__13959 (.I0(n10141), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), .O(n10142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__13959.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__13960 (.I0(n10140), .I1(n10139), .I2(n10131), .I3(n10142), 
            .O(n10143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__13960.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__13961 (.I0(n10134), .I1(n10137), .I2(n10133), .I3(n10143), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h01ff */ ;
    defparam LUT__13961.LUTMASK = 16'h01ff;
    EFX_LUT4 LUT__13962 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] ), .O(n10144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13962.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13963 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] ), .I2(n10144), 
            .O(n10145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__13963.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__13964 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] ), .O(n10146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13964.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13965 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] ), .O(n10147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13965.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13966 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] ), .O(n10148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__13966.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__13967 (.I0(n10145), .I1(n10146), .I2(n10147), .I3(n10148), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/qRVD )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__13967.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__13968 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13968.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13969 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13969.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13970 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13970.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13971 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(n10149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13971.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13972 (.I0(n10149), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13972.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13973 (.I0(n10149), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13973.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13974 (.I0(n10149), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__13974.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__13975 (.I0(n10135), .I1(n10149), .O(n10150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13975.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13976 (.I0(n10150), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__13976.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__13977 (.I0(n10150), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__13977.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__13978 (.I0(wVideoVd), .I1(\MVideoPostProcess/rVtgRstSel ), 
            .O(\MVideoPostProcess/qVtgRstCntCke )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13978.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13979 (.I0(\MVideoPostProcess/rVtgRstCnt[8] ), .I1(\MVideoPostProcess/rVtgRstCnt[9] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[10] ), .O(n10151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__13979.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__13980 (.I0(\MVideoPostProcess/rVtgRstCnt[4] ), .I1(\MVideoPostProcess/rVtgRstCnt[5] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[6] ), .I3(\MVideoPostProcess/rVtgRstCnt[7] ), 
            .O(n10152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__13980.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__13981 (.I0(\MVideoPostProcess/rVtgRstCnt[0] ), .I1(\MVideoPostProcess/rVtgRstCnt[1] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[2] ), .I3(\MVideoPostProcess/rVtgRstCnt[3] ), 
            .O(n10153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__13981.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__13982 (.I0(n10151), .I1(n10152), .I2(n10153), .O(\MVideoPostProcess/equal_18/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f7f */ ;
    defparam LUT__13982.LUTMASK = 16'h7f7f;
    EFX_LUT4 LUT__13983 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] ), 
            .O(n10154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__13983.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__13984 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[1] ), .O(n10155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__13984.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__13985 (.I0(n10154), .I1(n10155), .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), .O(n10156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13985.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13986 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_ack ), .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(n10157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13986.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13987 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[0] ), 
            .I1(n10156), .I2(n10157), .O(\MVideoPostProcess/inst_adv7511_config/n816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f1f */ ;
    defparam LUT__13987.LUTMASK = 16'h1f1f;
    EFX_LUT4 LUT__13988 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] ), .O(n10158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13988.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13989 (.I0(n10158), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] ), 
            .O(n10159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__13989.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__13990 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
            .I1(n10159), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] ), .O(n10160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__13990.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__13991 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .I1(pll_inst1_LOCKED), .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I3(rBRST), .O(n10161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__13991.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__13992 (.I0(n10160), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .I3(n10161), .O(\~ceg_net510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__13992.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__13993 (.I0(n10156), .I1(n10157), .O(n10162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__13993.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__13994 (.I0(n10162), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13994.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13995 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__13995.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__13996 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/n1107 ), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1235 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__13996.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__13997 (.I0(rBRST), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(ceg_net477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__13997.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__13998 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(ceg_net42)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__13998.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__13999 (.I0(\MVideoPostProcess/inst_adv7511_config/w_ack ), 
            .I1(n10156), .I2(ceg_net477), .I3(\~ceg_net510 ), .O(ceg_net1377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__13999.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__14000 (.I0(rBRST), .I1(\MVideoPostProcess/inst_adv7511_config/n1107 ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14000.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14001 (.I0(oAdv7511SclOe), .I1(iAdv7511Scl), .I2(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__14001.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__14002 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .O(n10164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14002.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14003 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n10165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14003.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14004 (.I0(n10163), .I1(n10164), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(n10165), .O(ceg_net567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__14004.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__14005 (.I0(ceg_net567), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(n10165), .O(n10166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__14005.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__14006 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n10167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14006.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14007 (.I0(n10163), .I1(n10166), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(n10167), .O(n10168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf10f */ ;
    defparam LUT__14007.LUTMASK = 16'hf10f;
    EFX_LUT4 LUT__14008 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(n10168), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14008.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14009 (.I0(n10164), .I1(n10167), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc102 */ ;
    defparam LUT__14009.LUTMASK = 16'hc102;
    EFX_LUT4 LUT__14010 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .O(n10169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14010.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14011 (.I0(n10169), .I1(n10167), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(ceg_net1421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h070c */ ;
    defparam LUT__14011.LUTMASK = 16'h070c;
    EFX_LUT4 LUT__14012 (.I0(n10167), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n10170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14012.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14013 (.I0(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_last_1P ), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__14013.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__14014 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] ), 
            .O(n10172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14014.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14015 (.I0(oAdv7511SdaOe), .I1(n10171), .I2(n10172), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcc35 */ ;
    defparam LUT__14015.LUTMASK = 16'hcc35;
    EFX_LUT4 LUT__14016 (.I0(oAdv7511SdaOe), .I1(n10173), .I2(n10164), 
            .O(n10174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__14016.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__14017 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n10175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14017.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14018 (.I0(iAdv7511Sda), .I1(oAdv7511SdaOe), .O(n10176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14018.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14019 (.I0(n10172), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .I2(n10176), .I3(n10164), .O(n10177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14019.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14020 (.I0(n10164), .I1(oAdv7511SdaOe), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14020.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14021 (.I0(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .O(n10179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__14021.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__14022 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14022.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14023 (.I0(n10179), .I1(n10180), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n10181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bb0 */ ;
    defparam LUT__14023.LUTMASK = 16'h0bb0;
    EFX_LUT4 LUT__14024 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .O(n10182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__14024.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__14025 (.I0(n10182), .I1(n10167), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14025.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14026 (.I0(n10177), .I1(n10178), .I2(n10181), .I3(n10183), 
            .O(n10184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__14026.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__14027 (.I0(n10174), .I1(n10175), .I2(n10184), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n10185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__14027.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__14028 (.I0(n10164), .I1(oAdv7511SdaOe), .I2(n10170), 
            .I3(n10185), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;
    defparam LUT__14028.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__14029 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I1(n10167), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .O(n10186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14029.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14030 (.I0(n10175), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14030.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14031 (.I0(n10164), .I1(ceg_net567), .I2(n10186), .I3(n10187), 
            .O(ceg_net1389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0dcc */ ;
    defparam LUT__14031.LUTMASK = 16'h0dcc;
    EFX_LUT4 LUT__14032 (.I0(n10175), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n10176), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .O(n10188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__14032.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__14033 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I1(n10180), .I2(n10167), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n10189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h50cf */ ;
    defparam LUT__14033.LUTMASK = 16'h50cf;
    EFX_LUT4 LUT__14034 (.I0(n10188), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I2(n10189), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__14034.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__14035 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14035.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14036 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n10190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14036.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14037 (.I0(n10165), .I1(n10167), .O(ceg_net617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__14037.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__14038 (.I0(n10164), .I1(n10172), .I2(n10175), .O(n10191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14038.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14039 (.I0(ceg_net617), .I1(n10190), .I2(n10166), .I3(n10191), 
            .O(ceg_net1460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__14039.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__14040 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), .I2(n10169), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__14040.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__14041 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n10193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14041.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14042 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n10193), .O(n10194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14042.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14043 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n10176), .I2(n10172), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n10195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__14043.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__14044 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n10196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfd40 */ ;
    defparam LUT__14044.LUTMASK = 16'hfd40;
    EFX_LUT4 LUT__14045 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] ), 
            .I1(n10195), .I2(n10165), .I3(n10196), .O(n10197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__14045.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__14046 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] ), 
            .I1(n10192), .I2(n10194), .I3(n10197), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__14046.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__14047 (.I0(n10165), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n10198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14047.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14048 (.I0(n10164), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I3(n10190), .O(n10199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1700 */ ;
    defparam LUT__14048.LUTMASK = 16'h1700;
    EFX_LUT4 LUT__14049 (.I0(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I1(n10169), .I2(n10198), .I3(n10199), .O(ceg_net1523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__14049.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__14052 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n10172), .I2(n10164), .O(n10201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14052.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14055 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), .I2(n10164), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__14055.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__14056 (.I0(n10180), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(n10201), .I3(n10203), .O(n10204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__14056.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__14057 (.I0(n10172), .I1(n10176), .I2(n10164), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__14057.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__14058 (.I0(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(n10180), .I3(n10165), .O(n10206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__14058.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__14059 (.I0(n10170), .I1(n10164), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(n10206), .O(n10207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d7 */ ;
    defparam LUT__14059.LUTMASK = 16'h00d7;
    EFX_LUT4 LUT__14060 (.I0(n10205), .I1(n10204), .I2(n10193), .I3(n10207), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff */ ;
    defparam LUT__14060.LUTMASK = 16'h10ff;
    EFX_LUT4 LUT__14061 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n10163), .I2(n10164), .I3(n10165), .O(ceg_net1531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__14061.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__14062 (.I0(n10165), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(n10205), .I3(ceg_net1531), .O(ceg_net1415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80 */ ;
    defparam LUT__14062.LUTMASK = 16'hff80;
    EFX_LUT4 LUT__14063 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n10193), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__14063.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__14064 (.I0(n10164), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n10208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14064.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14065 (.I0(n10169), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n10209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14065.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14066 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .O(n10210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__14066.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__14067 (.I0(n10209), .I1(n10208), .I2(n10210), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__14067.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__14068 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(n10168), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14068.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14069 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(n10168), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__14069.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__14070 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] ), 
            .O(n10211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14070.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14071 (.I0(n10168), .I1(n10211), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14071.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14072 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] ), 
            .O(n10212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14072.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14073 (.I0(n10212), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(n10168), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14073.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14074 (.I0(n10212), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I3(n10168), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__14074.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__14075 (.I0(n10212), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] ), 
            .O(n10213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14075.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14076 (.I0(n10168), .I1(n10213), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14076.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14077 (.I0(n10212), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] ), 
            .O(n10214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14077.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14078 (.I0(n10214), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I2(n10168), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14078.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14092 (.I0(n10164), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .O(n10220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14092.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14093 (.I0(n10220), .I1(n10167), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc102 */ ;
    defparam LUT__14093.LUTMASK = 16'hc102;
    EFX_LUT4 LUT__14094 (.I0(n10220), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .O(n10221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14094.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14095 (.I0(n10221), .I1(n10167), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc102 */ ;
    defparam LUT__14095.LUTMASK = 16'hc102;
    EFX_LUT4 LUT__14096 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14096.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14097 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14097.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14098 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14098.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14099 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14099.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14100 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14100.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14101 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14101.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14102 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14102.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14103 (.I0(n10209), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[3] ), 
            .O(n10222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14103.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14104 (.I0(n10209), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] ), 
            .I3(n10195), .O(n10223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__14104.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__14105 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n10224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__14105.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__14106 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I2(n10192), .I3(n10194), .O(n10225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14106.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14107 (.I0(n10224), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .I2(n10225), .O(n10226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14107.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14108 (.I0(n10222), .I1(n10223), .I2(n10165), .I3(n10226), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0ff */ ;
    defparam LUT__14108.LUTMASK = 16'hb0ff;
    EFX_LUT4 LUT__14109 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .I2(n10192), .I3(n10194), .O(n10227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14109.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14110 (.I0(n10209), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] ), 
            .I3(n10195), .O(n10228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__14110.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__14111 (.I0(n10228), .I1(n10165), .I2(n10224), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .O(n10229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__14111.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__14112 (.I0(n10227), .I1(n10229), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14112.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14113 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .I2(n10192), .I3(n10194), .O(n10230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14113.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14114 (.I0(n10209), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] ), 
            .I3(n10195), .O(n10231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__14114.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__14115 (.I0(n10231), .I1(n10165), .I2(n10224), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .O(n10232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__14115.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__14116 (.I0(n10230), .I1(n10232), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14116.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14117 (.I0(n10209), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] ), 
            .I3(n10195), .O(n10233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__14117.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__14118 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .I2(n10192), .I3(n10194), .O(n10234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14118.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14119 (.I0(n10224), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .I2(n10234), .O(n10235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14119.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14120 (.I0(n10222), .I1(n10233), .I2(n10165), .I3(n10235), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0ff */ ;
    defparam LUT__14120.LUTMASK = 16'hb0ff;
    EFX_LUT4 LUT__14121 (.I0(n10209), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] ), 
            .I3(n10195), .O(n10236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__14121.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__14122 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .I2(n10192), .I3(n10194), .O(n10237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14122.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14123 (.I0(n10222), .I1(n10236), .I2(n10165), .I3(n10237), 
            .O(n10238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__14123.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__14124 (.I0(n10224), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .I2(n10238), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__14124.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__14125 (.I0(n10209), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] ), 
            .I3(n10195), .O(n10239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__14125.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__14126 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .I2(n10192), .I3(n10194), .O(n10240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14126.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14127 (.I0(n10224), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .I2(n10240), .O(n10241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__14127.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__14128 (.I0(n10222), .I1(n10239), .I2(n10165), .I3(n10241), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0ff */ ;
    defparam LUT__14128.LUTMASK = 16'hb0ff;
    EFX_LUT4 LUT__14129 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .I2(n10192), .I3(n10194), .O(n10242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__14129.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__14130 (.I0(n10209), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] ), 
            .I3(n10195), .O(n10243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__14130.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__14131 (.I0(n10243), .I1(n10165), .I2(n10224), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .O(n10244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__14131.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__14132 (.I0(n10242), .I1(n10244), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14132.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14140 (.I0(oAdv7511SdaOe), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(iAdv7511Sda), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n10245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3 */ ;
    defparam LUT__14140.LUTMASK = 16'hedf3;
    EFX_LUT4 LUT__14141 (.I0(n10245), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n10246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14141.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14142 (.I0(n10208), .I1(n10175), .I2(n10246), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__14142.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__14143 (.I0(n10176), .I1(n10192), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n10247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0cd */ ;
    defparam LUT__14143.LUTMASK = 16'hf0cd;
    EFX_LUT4 LUT__14144 (.I0(iAdv7511Sda), .I1(n10198), .I2(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .O(n10248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__14144.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__14145 (.I0(n10164), .I1(n10247), .I2(n10193), .I3(n10248), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff70 */ ;
    defparam LUT__14145.LUTMASK = 16'hff70;
    EFX_LUT4 LUT__14146 (.I0(n10192), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(n10193), .I3(n10208), .O(n10249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__14146.LUTMASK = 16'he000;
    EFX_LUT4 LUT__14147 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I2(n10198), .I3(n10249), .O(n10250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__14147.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__14148 (.I0(n10164), .I1(n10170), .I2(n10250), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__14148.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__14149 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[1] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), .O(n10251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14149.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14150 (.I0(n10251), .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), 
            .O(n10252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14150.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14151 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), .O(n10253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__14151.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__14152 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[7] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[8] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[9] ), 
            .O(n10254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__14152.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__14153 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I3(n10254), .O(n10255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__14153.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__14154 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .I1(n10252), .I2(n10253), .I3(n10255), .O(\MVideoPostProcess/mVideoTimingGen/qVrange )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__14154.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__14155 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14155.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14156 (.I0(n10162), .I1(n10161), .O(ceg_net941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14156.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14157 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14157.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14158 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[1] ), .O(n10256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14158.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14159 (.I0(n10256), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14159.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14160 (.I0(n10256), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__14160.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__14161 (.I0(n10256), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), .O(n10257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14161.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14162 (.I0(n10257), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14162.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14163 (.I0(n10257), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), 
            .O(n10258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14163.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14164 (.I0(n10258), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14164.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14165 (.I0(n10258), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__14165.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__14166 (.I0(n10258), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), .O(n10259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14166.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14167 (.I0(n10259), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14167.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14168 (.I0(n10258), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), 
            .O(n10260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14168.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14169 (.I0(n10260), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__14169.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__14170 (.I0(n10260), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__14170.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__14171 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14171.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14172 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] ), 
            .O(n10261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14172.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14173 (.I0(n10261), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14173.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14174 (.I0(n10261), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14174.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14175 (.I0(n10261), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14175.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14176 (.I0(n10261), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] ), 
            .O(n10262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14176.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14177 (.I0(n10262), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14177.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14178 (.I0(n10262), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14178.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14179 (.I0(n10262), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14179.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14180 (.I0(n10262), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] ), 
            .O(n10263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14180.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14181 (.I0(n10263), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14181.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14182 (.I0(n10263), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14182.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14183 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] ), 
            .O(n10264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14183.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14184 (.I0(n10263), .I1(n10264), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14184.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14185 (.I0(n10263), .I1(n10264), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14185.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14186 (.I0(n10263), .I1(n10264), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] ), 
            .O(n10265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14186.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14187 (.I0(n10265), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14187.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14188 (.I0(n10265), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14188.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14189 (.I0(n10265), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14189.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14190 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] ), 
            .O(n10266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14190.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14191 (.I0(n10265), .I1(n10266), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14191.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14192 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .O(\MVideoPostProcess/inst_adv7511_config/n780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14192.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14193 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14193.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14194 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] ), .O(\MVideoPostProcess/inst_adv7511_config/n790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14194.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14195 (.I0(n10158), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14195.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14196 (.I0(n10158), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .O(\MVideoPostProcess/inst_adv7511_config/n800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14196.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14197 (.I0(n10158), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14197.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14198 (.I0(n10159), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14198.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14199 (.I0(n10255), .I1(n10252), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .O(n10267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14199.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14200 (.I0(n10267), .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), 
            .O(\MVideoPostProcess/mVideoTimingGen/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14200.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14201 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), .O(n10268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__14201.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__14202 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), .I2(n10268), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), .O(n10269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14202.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14203 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[1] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .O(n9980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14203.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14204 (.I0(n10269), .I1(n9980), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), .O(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__14204.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__14205 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .I3(n10254), .O(n10270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__14205.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__14206 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), .O(n10271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14206.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14207 (.I0(n10271), .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), .O(n10272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__14207.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__14208 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), 
            .I1(n10270), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I3(n10272), .O(\MVideoPostProcess/mVideoTimingGen/qVde )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__14208.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__14209 (.I0(\MVideoPostProcess/rVtgRST[2] ), .I1(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
            .O(\MVideoPostProcess/mVideoTimingGen/n267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__14209.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__14210 (.I0(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 ), .O(\MVideoPostProcess/mVideoTimingGen/rHSync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14210.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14211 (.I0(n10267), .I1(n441), .O(\MVideoPostProcess/mVideoTimingGen/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14211.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14212 (.I0(n10267), .I1(n3654), .O(\MVideoPostProcess/mVideoTimingGen/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14212.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14213 (.I0(n10267), .I1(n3648), .O(\MVideoPostProcess/mVideoTimingGen/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14213.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14214 (.I0(n10267), .I1(n3646), .O(\MVideoPostProcess/mVideoTimingGen/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14214.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14215 (.I0(n10267), .I1(n3638), .O(\MVideoPostProcess/mVideoTimingGen/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14215.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14216 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), .O(n10273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__14216.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__14217 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I3(n10269), .O(n10274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__14217.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__14218 (.I0(n10273), .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I2(n10271), .I3(n10274), .O(\MVideoPostProcess/mVideoTimingGen/qHrange )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80 */ ;
    defparam LUT__14218.LUTMASK = 16'hff80;
    EFX_LUT4 LUT__14219 (.I0(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 ), .O(\MVideoPostProcess/mVideoTimingGen/rVSync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14219.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14220 (.I0(\MVideoPostProcess/mVideoTimingGen/dff_41/i4_pre ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 ), .O(\MVideoPostProcess/mVideoTimingGen/rVde[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__14220.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__14221 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .O(n10275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14221.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14222 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14222.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14223 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14223.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14224 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n10278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14224.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14225 (.I0(n10277), .I1(n10278), .O(n10279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14225.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14226 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14226.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14227 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14227.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14228 (.I0(n10281), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I3(n10280), .O(n10282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100 */ ;
    defparam LUT__14228.LUTMASK = 16'h4100;
    EFX_LUT4 LUT__14229 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14229.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14230 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14230.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14231 (.I0(n10279), .I1(n10282), .I2(n10283), .I3(n10284), 
            .O(n10285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14231.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14232 (.I0(n10276), .I1(n10285), .I2(n10275), .I3(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__14232.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__14233 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .O(n10286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__14233.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__14234 (.I0(n10286), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .O(n10287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__14234.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__14235 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14235.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14236 (.I0(n10288), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .I3(n10277), .O(n10289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14236.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14237 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b */ ;
    defparam LUT__14237.LUTMASK = 16'hb00b;
    EFX_LUT4 LUT__14238 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14238.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14239 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I1(n10291), .I2(n10288), .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n10292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde */ ;
    defparam LUT__14239.LUTMASK = 16'hbdde;
    EFX_LUT4 LUT__14240 (.I0(n10290), .I1(n10292), .I2(n10289), .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n10293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__14240.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__14241 (.I0(n10279), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .O(n10294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__14241.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__14242 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b */ ;
    defparam LUT__14242.LUTMASK = 16'hb00b;
    EFX_LUT4 LUT__14243 (.I0(n10288), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14243.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14244 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14244.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14245 (.I0(n10295), .I1(n10280), .I2(n10296), .I3(n10297), 
            .O(n10298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccc */ ;
    defparam LUT__14245.LUTMASK = 16'h5ccc;
    EFX_LUT4 LUT__14246 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14246.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14247 (.I0(n10299), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I3(n10281), .O(n10300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcfa2 */ ;
    defparam LUT__14247.LUTMASK = 16'hcfa2;
    EFX_LUT4 LUT__14248 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bb0 */ ;
    defparam LUT__14248.LUTMASK = 16'h0bb0;
    EFX_LUT4 LUT__14249 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bb0 */ ;
    defparam LUT__14249.LUTMASK = 16'h0bb0;
    EFX_LUT4 LUT__14250 (.I0(n10299), .I1(n10283), .I2(n10301), .I3(n10302), 
            .O(n10303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__14250.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__14251 (.I0(n10300), .I1(n10303), .O(n10304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__14251.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__14252 (.I0(n10293), .I1(n10294), .I2(n10298), .I3(n10304), 
            .O(n10305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14252.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14253 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(n10280), .O(n10306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__14253.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__14254 (.I0(n10306), .I1(n10277), .I2(n10287), .I3(n10296), 
            .O(n10307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__14254.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__14255 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14255.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14256 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I3(n10308), .O(n10309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8af3 */ ;
    defparam LUT__14256.LUTMASK = 16'h8af3;
    EFX_LUT4 LUT__14257 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bb0 */ ;
    defparam LUT__14257.LUTMASK = 16'h0bb0;
    EFX_LUT4 LUT__14258 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14258.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14259 (.I0(n10310), .I1(n10281), .I2(n10311), .O(n10312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__14259.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__14260 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bb0 */ ;
    defparam LUT__14260.LUTMASK = 16'h0bb0;
    EFX_LUT4 LUT__14261 (.I0(n10309), .I1(n10302), .I2(n10312), .I3(n10313), 
            .O(n10314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14261.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14262 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14262.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14263 (.I0(n10288), .I1(n10315), .O(n10316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14263.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14264 (.I0(n10292), .I1(n10316), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1441 */ ;
    defparam LUT__14264.LUTMASK = 16'h1441;
    EFX_LUT4 LUT__14265 (.I0(n10307), .I1(n10314), .I2(n10317), .O(n10318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14265.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14266 (.I0(n10285), .I1(n10287), .I2(n10305), .I3(n10318), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__14266.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__14267 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14267.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14268 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14268.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14269 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14269.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14270 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n10319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14270.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14271 (.I0(n10319), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14271.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14272 (.I0(n10319), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14272.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14273 (.I0(n10319), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14273.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14274 (.I0(n10311), .I1(n10319), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14274.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14275 (.I0(n10288), .I1(n10319), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14275.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14276 (.I0(n10288), .I1(n10319), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__14276.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__14277 (.I0(n10296), .I1(n10319), .O(n10320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__14277.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__14278 (.I0(n10320), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14278.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14279 (.I0(n10320), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14279.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14280 (.I0(n10316), .I1(n10319), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__14280.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__14281 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14281.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14282 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14282.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14283 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14283.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14284 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14284.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14285 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14285.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14286 (.I0(n10322), .I1(n10323), .I2(n10324), .I3(n10325), 
            .O(n10326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14286.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14287 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14287.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14288 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(n10326), .I3(n10327), .O(n10328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14288.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14289 (.I0(n10328), .I1(n10321), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14289.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14290 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14290.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14291 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14291.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14292 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10329), .I3(n10330), .O(n10331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14292.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14293 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14293.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14294 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14294.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14295 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14295.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14296 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14296.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14297 (.I0(n10332), .I1(n10333), .I2(n10334), .I3(n10335), 
            .O(n10336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14297.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14298 (.I0(n10336), .I1(n10331), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14298.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14299 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14299.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14300 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14300.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14301 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10337), .I3(n10338), .O(n10339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14301.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14302 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14302.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14303 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14303.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14304 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14304.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14305 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14305.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14306 (.I0(n10340), .I1(n10341), .I2(n10342), .I3(n10343), 
            .O(n10344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14306.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14307 (.I0(n10344), .I1(n10339), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14307.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14308 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14308.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14309 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14309.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14310 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10345), .I3(n10346), .O(n10347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14310.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14311 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14311.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14312 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14312.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14313 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14313.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14314 (.I0(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14314.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14315 (.I0(n10348), .I1(n10349), .I2(n10350), .I3(n10351), 
            .O(n10352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14315.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14316 (.I0(n10352), .I1(n10347), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[4].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14316.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14317 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14317.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14318 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14318.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14319 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14319.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14320 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n10356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14320.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14321 (.I0(n10353), .I1(n10354), .I2(n10355), .I3(n10356), 
            .O(n10357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__14321.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__14322 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14322.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14323 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14323.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14324 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14324.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14325 (.I0(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/rWA[0] ), 
            .I2(n10359), .I3(n10360), .O(n10361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14325.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14326 (.I0(n10358), .I1(n10361), .I2(n10357), .I3(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[5].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__14326.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__14327 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14327.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14328 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14328.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14329 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14329.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14330 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14330.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14331 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14331.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14332 (.I0(n10363), .I1(n10364), .I2(n10365), .I3(n10366), 
            .O(n10367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14332.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14333 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14333.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14334 (.I0(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(n10367), .I3(n10368), .O(n10369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14334.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14335 (.I0(n10369), .I1(n10362), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[6].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14335.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14336 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[1] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .O(n10370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14336.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14337 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14337.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14338 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(n10370), .I3(n10371), .O(n10372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14338.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14339 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14339.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14340 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14340.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14341 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14341.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14342 (.I0(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14342.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14343 (.I0(n10373), .I1(n10374), .I2(n10375), .I3(n10376), 
            .O(n10377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14343.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14344 (.I0(n10377), .I1(n10372), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[7].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14344.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14345 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14345.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14346 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14346.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14347 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10378), .I3(n10379), .O(n10380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14347.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14348 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14348.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14349 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14349.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14350 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14350.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14351 (.I0(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14351.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14352 (.I0(n10381), .I1(n10382), .I2(n10383), .I3(n10384), 
            .O(n10385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14352.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14353 (.I0(n10385), .I1(n10380), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[8].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14353.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14354 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[3] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n10386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14354.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14355 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14355.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14356 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[9] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14356.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14357 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14357.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14358 (.I0(n10386), .I1(n10387), .I2(n10388), .I3(n10389), 
            .O(n10390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14358.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14359 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14359.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14360 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14360.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14361 (.I0(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(n10392), .O(n10393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__14361.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__14362 (.I0(n10391), .I1(n10393), .I2(n10390), .I3(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[9].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__14362.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__14363 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14363.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14364 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14364.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14365 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14365.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14366 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[9] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14366.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14367 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14367.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14368 (.I0(n10395), .I1(n10396), .I2(n10397), .I3(n10398), 
            .O(n10399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14368.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14369 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14369.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14370 (.I0(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(n10399), .I3(n10400), .O(n10401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14370.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14371 (.I0(n10401), .I1(n10394), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[10].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14371.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14372 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n10402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14372.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14373 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14373.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14374 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(n10402), .I3(n10403), .O(n10404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14374.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14375 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14375.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14376 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n10406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14376.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14377 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14377.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14378 (.I0(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .I2(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14378.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14379 (.I0(n10405), .I1(n10406), .I2(n10407), .I3(n10408), 
            .O(n10409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14379.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14380 (.I0(n10409), .I1(n10404), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[11].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14380.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14381 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14381.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14382 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14382.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14383 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14383.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14384 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14384.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14385 (.I0(n10410), .I1(n10411), .I2(n10412), .I3(n10413), 
            .O(n10414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14385.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14386 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14386.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14387 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14387.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14388 (.I0(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14388.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14389 (.I0(n10417), .I1(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/rRA[7] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I3(n10416), .O(n10418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100 */ ;
    defparam LUT__14389.LUTMASK = 16'h4100;
    EFX_LUT4 LUT__14390 (.I0(n10415), .I1(n10418), .I2(n10414), .I3(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[12].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__14390.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__14391 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14391.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14392 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14392.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14393 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14393.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14394 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14394.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14395 (.I0(n10419), .I1(n10420), .I2(n10421), .I3(n10422), 
            .O(n10423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14395.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14396 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14396.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14397 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[11] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__14397.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__14398 (.I0(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14398.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14399 (.I0(n10426), .I1(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/rRA[7] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I3(n10425), .O(n10427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100 */ ;
    defparam LUT__14399.LUTMASK = 16'h4100;
    EFX_LUT4 LUT__14400 (.I0(n10424), .I1(n10427), .I2(n10423), .I3(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[13].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__14400.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__14401 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14401.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14402 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14402.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14403 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[3] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n10430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14403.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14404 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14404.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14405 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n10432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14405.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14406 (.I0(n10429), .I1(n10430), .I2(n10431), .I3(n10432), 
            .O(n10433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14406.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14407 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14407.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14408 (.I0(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(n10433), .I3(n10434), .O(n10435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14408.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14409 (.I0(n10435), .I1(n10428), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[14].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14409.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14410 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[12] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[12] ), 
            .O(n10436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14410.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14411 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n10437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14411.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14412 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n10438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14412.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14413 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(n10439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14413.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14414 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n10440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14414.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14415 (.I0(n10437), .I1(n10438), .I2(n10439), .I3(n10440), 
            .O(n10441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14415.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14416 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[11] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[11] ), 
            .O(n10442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__14416.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__14417 (.I0(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(n10441), .I3(n10442), .O(n10443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__14417.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__14418 (.I0(n10443), .I1(n10436), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[15].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__14418.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__14419 (.I0(\genblk1.genblk1[0].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[0].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__14419.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__14420 (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1] ), .I2(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[2] ), 
            .O(n9781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__14420.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__14421 (.I0(n9781), .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] ), 
            .I2(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] ), .I3(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] ), 
            .O(n10444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__14421.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__14422 (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] ), .I2(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] ), 
            .I3(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] ), .O(n10445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__14422.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__14423 (.I0(n10444), .I1(n10445), .I2(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] ), 
            .I3(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] ), .O(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__14423.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__14424 (.I0(\genblk1.genblk1[1].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[1].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[1].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[1].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__14424.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__14425 (.I0(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[1].mPulseGenerator/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14425.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14426 (.I0(\genblk1.genblk1[3].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[3].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[3].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__14426.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__14427 (.I0(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[3].mPulseGenerator/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14427.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14428 (.I0(\genblk1.genblk1[4].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[4].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[4].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__14428.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__14429 (.I0(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[4].mPulseGenerator/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14429.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__14430 (.I0(\la0_probe18[0] ), .I1(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneLs ), 
            .O(la0_probe10)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__14430.LUTMASK = 16'h6666;
    
endmodule

//
// Verific Verilog Description of module EFX_FF_0129fa4d_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_0129fa4d_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_0129fa4d_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__5_5_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__5_5_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__5_5_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__5_5_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__16_16_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_SRL8_0129fa4d_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__1_1_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_0129fa4d__8_8_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_0129fa4d_221
// module not written out since it is a black box. 
//

