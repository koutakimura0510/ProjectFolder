//----------------------------------------------------------
// Create 2022/4/20
// Author koutakimura
// -
// SPI 通信を行うモジュール
// 
//----------------------------------------------------------
module fmbWrapper (
    output      oCs,
    output      oSck,
    output      oMosi,
    input       iMiso,
    output      oWp,
    output      oHold,
    output      oData,
    input       iAddr,
    input       iCke,
    output      oVd
);




endmodule