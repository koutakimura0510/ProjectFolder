//----------------------------------------------------------
// KEY Bit値
//----------------------------------------------------------
localparam SW_B     = 0; //0x04
localparam SW_DOWN  = 1; //0x02
localparam SW_UP    = 2; //0x01
localparam SW_LEFT  = 3; //0x20
localparam SW_RIGHT = 4; //0x10
localparam SW_A     = 5; //0x08