//----------------------------------------------------------
// Create 2023/10/14
// Author koutakimura
// -
// HyperRam Port Unit
// 
// 
//----------------------------------------------------------
module RAMIfPortUnit #(
	parameter pRamAdrsWidth	= 19,
	parameter pRamDqWidth = 8
)(
	// SRAM I/F Port
	output	[pRamDqWidth-1:0] oSRAMD,
	input	[pRamDqWidth-1:0] iSRAMD,
	output	oSRAM_nRST,
	output	oSRAM_nCE,
	output	oSRAM_RWDS,
	output	oSRAM_pCLK,
	output	oSRAM_nCLK,
	// Common Port
	input	[pRamAdrsWidth-1:0] iAdrs,
	input	iCmd,  // "1" Read, "0" Write
	input	[pRamDqWidth-1:0] iWd,
	output	[pRamDqWidth-1:0] oRd,
	output	oRvd,
    // Clk Reset
	input	iRST,
	input	iCKE,
	input	iCLK
);


//-----------------------------------------------------------------------------
// 調停が必要ない場合 50Mhz で動作可能
// それ以上はタイミング調整のロジックが必要
// 
// 50Mhz で動作させた場合で CLK遷移で Setuo/HoldTime は確保できるため、
// ユーザー側で特別な制御をする必要がなくなる。
// そのため、アドレスや書き込みデータはスルー制御とすることができる。
// 
//-----------------------------------------------------------------------------
reg  [pRamAdrsWidth-1:0] rAdrs;
reg  [pRamDqWidth-1:0] rWd;
reg  rOE, rWE, rCE;
wire [pRamDqWidth-1:0] wRd;
reg  [pRamDqWidth-1:0] rRd;
reg  rRvd;

always @(posedge iCLK)
begin
	rAdrs 	<= iAdrs;
	rWd 	<= iWd;

	if (iCKE)
	begin
		rOE <= ~iCmd;
		rWE <=  iCmd;
		rCE <=  1'b0;
	end
	else
	begin
		rOE <= 1'b1;
		rWE <= 1'b0;
		rCE <= 1'b1;
	end

	if (rWE) rRd <= iSRAMD;
	else  	 rRd <= rRd;

	if (iRST)		rRvd <= 1'b0;
	else if (rWE) 	rRvd <= 1'b1;
	else  			rRvd <= 1'b0;
end

assign oSRAMA = rAdrs;
assign oSRAMD = rWd;
// assign oSRAM_LB = 1'b0; // 常に有効
// assign oSRAM_UB = 1'b0; // 常に有効
// assign oSRAM_OE = rOE;
// assign oSRAM_WE = rWE;
// assign oSRAM_CE = rCE;
assign oSRAM_OE = 1'b1;
assign oSRAM_RWDS = 1'b1;
assign oSRAM_pCLK = 1'b1;
assign oSRAM_nCLK = 1'b1;
assign oSRAM_nCE = 1'b1;
assign oSRAM_nRST = 1'b1;
assign oRd = rRd;
assign oRvd = rRvd;

endmodule