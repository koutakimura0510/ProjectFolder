//////////////////////////////////////////////////////////////////////////////////////////
//           _____       
//          / _______    Copyright (C) 2013-2022 Efinix Inc. All rights reserved.
//         / /       \   
//        / /  ..    /   
//       / / .'     /    
//    __/ /.'      /     Description:
//   __   \       /      Top IP Module = efx_csi2_rx_top
//  /_/ /\ \_____/ /     
// ____/  \_______/      
//
// ***************************************************************************************
// Vesion  : 1.00
// Time    : Tue Aug  2 22:21:19 2022
// ***************************************************************************************
`define IP_UUID _rx
`define IP_NAME_CONCAT(a,b) a``b
`define IP_MODULE_NAME(name) `IP_NAME_CONCAT(name,`IP_UUID)

/*module efx_csi2_rx_top #(
    parameter HS_DATA_WIDTH = 16,
    parameter tINIT_NS = 100000,
	parameter CLOCK_FREQ_MHZ = 100,
    parameter NUM_DATA_LANE = 4,
    parameter PACK_TYPE = 4'b1111,
    parameter AREGISTER = 8,
    parameter ENABLE_VCX = 0,
	parameter FRAME_MODE = "GENERIC",    //1-ACCURATE, 0-GENERIC
    parameter ASYNC_STAGE = 2,
    parameter PIXEL_FIFO_DEPTH = 2048
)(
    input logic           reset_n,
    input logic           clk,				//100Mhz
    input logic           reset_byte_HS_n,
    input logic           clk_byte_HS,
    input logic           reset_pixel_n,
    input logic           clk_pixel,
    
    input   logic                       RxUlpsClkNot,
    input   logic                       RxUlpsActiveClkNot,
    input   logic [NUM_DATA_LANE-1:0]   RxClkEsc,      //
    input   logic [NUM_DATA_LANE-1:0]   RxErrEsc,
    input   logic [NUM_DATA_LANE-1:0]   RxErrControl,
    input   logic [NUM_DATA_LANE-1:0]   RxErrSotSyncHS,
    input   logic [NUM_DATA_LANE-1:0]   RxUlpsEsc, 
    input   logic [NUM_DATA_LANE-1:0]   RxUlpsActiveNot, 
    input   logic [NUM_DATA_LANE-1:0]   RxSkewCalHS, 
    input   logic [NUM_DATA_LANE-1:0]   RxStopState,   
    input   logic [NUM_DATA_LANE-1:0]   RxSyncHS,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS0,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS1,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS2,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS3,    
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS4,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS5,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS6,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS7,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS0,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS1,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS2,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS3,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS4,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS5,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS6,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS7,
    
    //AXI4-Lite Interface
    input                 axi_clk,
    input                 axi_reset_n,
    input          [5:0]  axi_awaddr,//Write Address. byte address.
    input                 axi_awvalid,//Write address valid.
    output logic          axi_awready,//Write address ready.
    input          [31:0] axi_wdata,//Write data bus.
    input                 axi_wvalid,//Write valid.
    output logic          axi_wready,//Write ready.
                          
    output logic          axi_bvalid,//Write response valid.
    input                 axi_bready,//Response ready.      
    input          [5:0]  axi_araddr,//Read address. byte address.
    input                 axi_arvalid,//Read address valid.
    output logic          axi_arready,//Read address ready.
    output logic   [31:0] axi_rdata,//Read data.
    output logic          axi_rvalid,//Read valid.
    input                 axi_rready,//Read ready.
	
    output logic          hsync_vc0,
    output logic          hsync_vc1,
    output logic          hsync_vc2,
    output logic          hsync_vc3,
    output logic          vsync_vc0,
    output logic          vsync_vc1,
    output logic          vsync_vc2,
    output logic          vsync_vc3,
    
    output logic          hsync_vc4,
    output logic          hsync_vc5,
    output logic          hsync_vc6,
    output logic          hsync_vc7,
    output logic          hsync_vc8,
    output logic          hsync_vc9,
    output logic          hsync_vc10,
    output logic          hsync_vc11,
    output logic          hsync_vc12,
    output logic          hsync_vc13,
    output logic          hsync_vc14,
    output logic          hsync_vc15,
    output logic          vsync_vc4,
    output logic          vsync_vc5,
    output logic          vsync_vc6,
    output logic          vsync_vc7,
    output logic          vsync_vc8,
    output logic          vsync_vc9,
    output logic          vsync_vc10,
    output logic          vsync_vc11,
    output logic          vsync_vc12,
    output logic          vsync_vc13,
    output logic          vsync_vc14,
    output logic          vsync_vc15,
    
    output logic [1:0]    vc,
    output logic [1:0]    vcx,
    output logic [15:0]   word_count,
    output logic [15:0]   shortpkt_data_field,
    output logic [5:0]    datatype,
    output logic [3:0]    pixel_per_clk,
    output logic [63:0]   pixel_data,
    output logic          pixel_data_valid,
    output logic          irq
);*/

`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
m0UtrF0XScYpp2IaD12i22iPkmzw4kq5Mtd3AQ01SgeZFZuwevsD8EOgOSl/J+fy
iJAVjrantkGGUNMWkl8F9vpvOjakXLqFZjz9BETriT/Gc/yj1VBKq8itcNGMPNNh
FySRgVPFVJT1vVG1tsqRv5ZKzJd5Zteu0fGZxUw3Xy9q2HF/PCI22X98YmgQuhGG
F4p+0Oe/iKNkfLBfP/XNbDOkw9RJ87SHY31Lun85/Zew7/zmqIvJFtfA8as8w3ix
lHkkKWKNb6pU8TpLl8MuMoZYkNaE64QL9iz0GGlGXZ7oo3R/BuXCyk2hl4dY8tj4
Bb54KZ/Hph2TjleedhU08Q==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 944 )
`pragma protect data_block
n+X6vee00jYnUz9BU/UXcT2HebHuUCu33lvDoGWCMG0DmG4O6gHfNnWUHwSUxzsc
ei+ED9sX8ybEfMQ9lzTx6tc/dK6//6cogQA9M9U+swHkQBwlk1NT+E/sSP9Cat2D
lh7hlZ9hxtMoEjtaay/0JVLURSJnjTqhx2kmW0VAqhbiyryzEMJbiQspdvzdiJy3
viiWSLSHGk4m5m529rzyuYSVm1wtq5TIhlEZNUVgN03DTfDBh8QzodFbzAb9Djhx
dwQKDBNKqv8OJd/ZNPzCYc0w9xgAM95j9ho3TZQeGi51JB8eA5vshXQMi4MAkLfB
DfTGyZaUElb0a5URY0SHDXWxWCRh/trlQZMOPN1ZIUC2hundlrJOtR5pJjHMc7mD
P3dB2FceU3mHwD1bGVFWLUV/gKjFW28YAi+jKrlwZpZU40X8/NGtkUgvlKhVq02G
KuPUr0hYwnJuljsWZyhSggGI6eS8JuPKfl21bY+RKLiJNU87n/JEDpy2/zrUKEz3
WH07o4S/2hhgPon1KoE3bMq1fVLRsSJCOFQuBBlf41SYICqAyv3qA/E6ztOb+O4r
KLXbM27kNlTqum5RPXjiKacTRG1MuLbOkiuBHA+Z79NSA0gwKFa6NjSGZ6N7AFj7
113OSOQMlz7mH4k7V6d+sdcd8c9Uzld20PcxCkq9d79KF3fPB8tPRDuRvXUT1jXF
66w5JhdXZDfaPolet3BUTlyTmEkORZPgnYLq8vNqx+GUxR22YTRRuSyTYUE2S0in
jWRiv9V9srd3qbFqyw/f16Rxr3+SkG8GeVFbox1eqvrS+QWkHtztr4BjEptk1UPB
A48v5Tl1K3SF/bxrGRos5+OzwK+gio2XDG+bZ9r5Ouu6DK154Dal4YOMQQesJXRI
BhAbJSqOsYNW0gk1WDM821yzUhN32fOz1aamlCHTzbUdkFo3Whakgi28ciY11bP1
WEh3aWxLjgufCEFKXvyKpZl/TjrZbP/OnsBEM61f25PPhVGGU+7R0I3fZOe1KKvQ
Urf1uuycLyh5H/cbWvVlEuX4Yo4kU4aux3yP+do2OaUB5CEO7NvACp/3Qhe89K2U
OBpBy7y5U9tuCNy7xKcfRvEBOFvt85Y8/NV1TiP1Qa9SYaT6UCHXXyUPsMOiQmyk
hsecMf54Do64G1XZLHvDLCukXCOhAFTxf5hex4PYxkuVFhZMMMYZXVx/LzUjQ/+y
8tUSbutoYb6eHIiC5cOGvwVg7arVxCCAauhwBLS6zp4=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
guG1hKDQP5Iof2xzDc/03pYHi8KTUjFe/Q+P9DrCmdBQE4z+YUaLDYCt+UkCk2P2
UybtnfhF92svVVknwh9qd9AUdGiDGwbGsLXqBQRQCGuqC3wWWbVi3VrGrY8FzvnN
yuZJMrTLuaSCHmcODrjYnLWHRuh7Oa5t7EJvivvAIUz7fCr1oFeHrvwselSUlE8i
Lgm7Bp3AwY6roAV5sS8RopZ0MLHgysf4PiPHK6lImUmlbWvsaQ4O+TXtvMzfsZXI
+2O/urs4i5RFvxye5DCG093uBces2QTaTwPQDDRlJqHrwYAopoLg7a8a4Fj7YH+e
mg1HNFVyr5wiOOHq48SAZA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 25408 )
`pragma protect data_block
SVytidGo/9tkIfiS6YpbEcNFZSQoQR1llCjDRUCmIli5152sTUyhgWsyyiw9ooQy
is1sCW3NNRo24P6QrsY5Zwz2XdZF/W98H9Xl97kevFXMmxoV38bcBy096N+PW9oA
2HBhb11fO16LMuM0Zp6TkGXr5YfLOST1nzBVpZnCJGE4US8+wL7zdbDq2MbIPxOz
QQ7rhSrsqmkjG0DojlYtP5/ZJoke1sZJ+K8OokESnN8yggFZZj+kYOcBmMYERBNH
Y4PInF7YTN1xrZh7wi1cz+wemIEGV52ypNdQQS0wjUKxbG0NQVWL2yPKV1FtFWh8
c57JUNUpMjlSHeM+dZN9t2EPw8Z0TjtdvmYjZtqlcWldTa2+Wxkwp9Z1XYfhWLLM
MRAdZkCetB5Oe1OYAkPIdZIWd3kMkH5CiBc9MCcXDHe9x4eblcXONHKEgaqR557a
xiacNPCFwMfZEHsHSO45i73tKTQOQtm0I2419GPT0hxA5VhE8JbJh9Lg7LbjFKRB
JlGydKHyDyK1DhsTgZyYy46rjgG0F+WWj/ipkHJXxRkKPEKC4LrS0XeI7GmaQjZO
Z/5si0eU4MLG0MrXwockVoWyAavKVgIPPV9U0mPxbgWhMFHEf9egBywCNCFvAFpM
rQKXKCOr4MezhgJ9UCNal4d3vnrqD9aKHuc+SX5AgiMCwp+/mg0/cOdvZ+TppDHb
L+KYAgqEt+kLWl2qsKU7rXBa5av0wnjqfo15nmYGxLw7vI/W9yffaH5frD/JiQne
9Gm8Kkm1sMeU86dsHjOr98GYoCNb8GVG4WaPH9W7jRVd66Mpy88NjAUNnDAVmvqn
MRdllu/LgLRxSVOGE35pc811vrV1/ZZUXHSc6/H4aR2107KIAo8yOw4l5OUEIgj8
HMMXbVW5is3pmrGz+NxVfcgBFtWf4I6EWUeTPCb8/sg8LnSP3+4f5pPebVG5mKOm
5GzekEFE0Zd8XcdNhYoKRP9ninB3fOjm7XWR04G0zShbV+f9R1HyLcSqCAh2xVt2
veZQ7DWGFiNl1tif2ARc5zgLoOPwMNxAz5hP7GlcQZLF1w+rri4k2/1xLtf5bQAh
T51MI6Q8D4NFIAYNOhk6R+XD8sidvDSaQzkvfnFW00h2HHzjt9cQS9YPxqRHBAn4
4w0deM0MAaRRb39x2ilAFW8zaNryxJLk4hnu9pSoUk1v5XYaPdQwy6DL62Upu/7z
hz6ZZPaaZjyd0VY8DQBpv2n0oxuIdH1cDdvwjlRhaU0RbVfPsimDLJwdNeRGS2BR
Yvh9OUuQNZmvuy3TU/ptG7TpHqD62hFaxTUvfNBJqDyWsE7rgL5Fh7Tox6b61OFC
ASGAXdVezcWjnVwYuZ4dSGHTpKZ58svdfvdHLis9mXVq//LImXNdBuLz8ez838Rt
MpjCHPoOZ83vOCOfJCA1zgTkrP5yhtP7SDoQFtaLk+BT2bnXhUC/Vuj6/wIg1ZaL
kqF2vG7lJivzs3O1ckR8dlLR4VDtLSJyr0edkbp8SIcNvsnA6c9iFXaK7YLOtOcA
PETF75s+VyKsw6MjMDq6aPNaaU1dAbvMdtuPcDDhulHU1brUOA/W2uhCpUsaDYzU
G0hDbGFMB/f8YA1vMbOUQ0UEZvDuM6RgBEuw0nem1CamG6QikqiL7y0ismZVn0AR
JloiTB+G08BeF2NzctHyWDQP7ysCdgV3Cj9ZpRwiAcrg4XUlZq47p4Oe+pu7MAXi
z5JBZ9KkBr9FZSyjomZAOiAbIJk2r3RhA9tIgmVj4dHCVcVeo/uKNLlbTSPErnql
gBbLPiH/nLy57wL/iOOFB/h9D+XjlOnLSsOmOvV/Ge1bI7qtK4XWQYxTMbQFBDtJ
Spb/HLnukLOyzJJ8DxtNbsSYDz/XD1bFZHuvDh/AHLrMQi/Jb1X2bwONj4ZcA/U5
qIpbLry1N20t3dc6/UJS7cEaNrVoBGW+Gc98jBtBj/HpzoXAwk7ossdibj3FcVOW
P5ycdDYCUCfUk8UipNWibioK39Kywl0t4LZ67FCj3j6/sLg2YQ+xIpjDQMWqx5BY
5ANGiAFFGp1w+Snmp2JPQ3F3Z9EBgiLDoualZLwScTvZ1Rrivlfiah7LNofKGp52
ckJhkFcI0KTRX/hm2SG8ekW9HGr4im/4ONJvOIGAt77GyQ/+FLb1QTTOs0kp6b9o
YR+679nf5LbbiHS/UnxqR88jmacsm3F3nnl/kuZhs4hyMvE04s73TxK3d4C1FXL1
7xYEFZc1kQk8RYKk4wbGD0g9dpc/Ed0kAyiiF0qn8YqCRgkzp4ev70Hp2EKVb9/J
oivIleQn51fZrpJGWYJxoMHWQyy1/uwDreLPrFqBlbWjxCuFp+p3eC/0RZiXz3sU
ka5RELBSIZiFpjpUFiQw6OgNnEKmcFKbdo1mcaHkUVIct2klxXTQXBH0/eNFIDZU
XfyZqRq2Gi+dGgQ7llyIhn6E1dOpEkqGgGoj9TKlSpMiinX7YF7/YWRIgwSoTpf5
VO+C6LHW0aP0h8xJ92A3f3hRkosY+jlaHUphjv/vy9bGrMGtYW65Ox0cQMxYgXvf
YcNfNS9NpADt7cgyI8wTDbY9uvfN+ggQ4iFbza3ejW0FG7GDKWtMwmzCahMgDqaI
LtXOyxxqtoVvsL/FZX30cq3R6b0nCu08wtSPfFDJntd9odeb7oiFmZ/DblNFEty8
9kdyqwLHL0MpnIZe36jws6hOOHXu7m3efiTgtYE5ARyKWaQvKq97W/MOT5VTmlrN
gJl0PldQfcrYn98bTGwt4lTgJ7n+uyNW/tXsK3mq28DrCCU+iEbi4crJbAEMXulb
Mj0GhrZsuEf40UVLj06wQPrNfc4YPxVoLoQRZFBDqMi5/1yaEI2JNTgHRxz9gj7I
UjYg4uLEk8wCUzgOpdiNvtIHsbpVN+qbpFSFr+XELwZ2uRIcumLh4NopwNTWWDFr
6WKqqpi1GabxtNjJxeoQNe6WLZyeB7MfD5IZcLuc5NY1jeMkfjxrAoGvL9qDjnaT
j6aP5nptqFnzjyg4Hp+znSMphN9XrE/F2lt/OHJCN3Xw9fHJv8U4TyRcnn4Tf/GE
e6ml4tE8TOr6UDWr6FybUe75J8h5V4dPX1G+waZfyBLt7Cne0TI/EQ5AJdqCb3bo
ELSUa4XXjb1WuPdBniHxIyjEQKYW9SNm7pdR46RFyOHdp+bbwO3UWdsw0Yx4v91O
oVarEA4jtZPyBNxO78wkMegIxyyio9coN1I12o03koF9MeYgvzHaUERTTrYarOz7
UUcJBA32nyJLvITZKGNAafjmTzjt6ZsZsL2baiS99QrI8Fh95mG29e/t0mw+Vwr2
7X9aygUDWLD185skPoAjFdJyeBRcp9n1I75OoBetays580fj8mTXx6ApvyFr8u5P
PhXZTvjb0vlvFrohqV7ywxPS3N1rPoP6C4uwoDMOI9tb6crl9M274A8O8WEKoANp
fkqH43V85ScVT+bvJfDvj373djWbDxPbCFcTAPRbPDf9kSva+8274BZegOIe5L2z
ZqElBEo9+dShARjUWrhCC9JdQr7J5R7saDmY9cD8AuIVx0WK2dMp7ktJsvJ+e4ag
FGmGuGrO6NsONOHVttIMMoE+fh4VCqLuGYq1hKTKTs8o96S3VtLuckp1/E66hR5x
rK9VkMVBDZpSJVCokBPwWB/oVTcasnDa8DqkAkf/s7acZ7DtspGxUsolKflOhDo4
o47sKQywBFmKqejjmM78f7qGmaonFI/BYsUl+Oc7jVXiSHkYEY7vjjalbtPwaUor
62hPKqxJPTICXm/gwBDJqefnOiffoufpF4NzuaD3Z3z72tv+HZZFd6xW6Xg1wTlh
JzrehVS2YxkHdDa7SfXkXFJwxXNDHf4FOp3sfCUxpwS5SWJ5OiY8KTZt7LDDh0U/
KRG/UDsL/czs9+AMHu0ge/TEKEHbS+cI4+FtiG0zs8vQHk+hF02SVNtgISQvV55r
I5S2VadiPbX+orlqE38yWaQvf1WeeO7eSCTy2m3K6tE38rT2TeeT+Iuc6iVv4Rr0
xOswFHPVYYJiqmTG0LN7YQTZ36VIBLxD58PqcSm+0Vg17ryACdXbyH5ZOuZzR43z
ubSVvDwgmLyXmvswRukwnfWUPoPW+YRjzP5110SCEnwxnjCvLKPFVM5Gw6OyDpaQ
fw8KPG9QhFZKLkv3pQ6BfaO2Ss9WLSPU2ZIMgJawBO9Ke5KRH1mUIzyB1GJ/qQnj
0+T93fwcDWKYYqDeSt63fK3VdmgHANAlj7qQidva3XdR4Ww1PgkMXyBSPptAZXJ5
YvUrnY/q3qcyb7Uf39eZFvn3imyrCp5rGg/VmQLgNNw+M6mN8JjUgco7UOz5arLz
BP9B24QyxcmoPiho4VgeLr0tookGLYg3N++6SFV25AbA/OQqDC5ys5oCV+Sy5eQT
SYzsspUBt4RB4M9RpkkuCdtgjhRVa9WAhfSnuxGrRic2t7lPORsWOAOvdmpGO9YH
Y40+BIl0jLUrfyWCBT2KCKNVk/RKDxybxfn8H0gNWCjzc6JZWPKv1P1aGQNWbMrd
AyJ8dkq8Qy7im6b59EJ62Jksr/XB5mH6yv1FmGNnKigethOkB2/gc+yPngG07Mfe
SlhdDoPy+qB+U+nLS8yC4op77rdcsUU6exwZWvnSDVOyaqhfNvMYobUT7iOEY4se
Fx+h/sGIeX8nzDL5cm0qPE0AxPDy6dsrsrq95obbRuvRWjtuU4ax/gWhJUtYkLWF
33pWtwAXbElbNMGc45Z4K6dlQTq1wqLvE8ZWfxkK/tNFmEfOhp56nUuTjYdNOtPN
hm19NNjJS+Q9OHeMpHu3qEQY3m4iyZ/zkOZkDLzjH5VN6ni+YaOBp7wFy61EjEWs
Uy4EdSzeDDajkyXHV914G0W/4dSYW7ZWz5I7Gz+/Qrl7RBKwCsA+IZMU19NEW+zU
o5CEnBuo1gFZNJRhQOQVVlv0+LN+Q07QZSVD9OgrTo0sHq6XAyJ0l/e7FlqtGw3B
WfSobj+zA0TVRjOFTf2uhirzPn8AQSUrrcgWF1WwlqiTFJSbuaTlKwzee9NDqt8P
Nu+3Ejt9+ms7m4CZsUROFxWeWv7P/l3a9i9OnOMe0ulWatWdpDlFyNVuUYDuxb5P
xUypV3tcFYR2ub4ezaQF/bIetxNil++e//HdicOJ6BQ43lisoLOfSnKn7kXf27aE
BdXiSWYp08SJCZSKp3gAPnB2wVkG9GhvI7gcm8JAhOEOk5XK1Zh1pNNiIDyX7s99
IMsZah8iUQHvCxlatulZPLuPOp36+LpOjLKtydTJhHNQ9YE9qWDqpLSMnZA9L9KM
TH7aXnXZ98nQpKO0a2V+SfU65flYtvMK0L0mhT7KNLyyxrwyIWEIuQwVxuYSbk2e
/iqemBVBKKbd+4oMSrJ0OuQwGiL7xODONXgEkF7xm3l44tfsowRKhQVFEQ5B3Us3
AuZtOfr780IxXm6/jU0q66TI2CLOHTUEQetq4WOrAmc4wQSeSQmR4rKaRtMtPD+Z
xV/jGIJ8wH5QrP6D3I5dsOrlgaM/50WGfR5vgC0/xn34dTIAg4e8prSHGRlhw+g1
pyLZzWlpHjxtfCHDRPR9v0VVLRDbO2NDQQeU0Gh4SUXQ9aoTEmSf1GCG48dP1kA7
CKQAsxtC8u4lOyHyuhKoww7so8RMjH3100naQOyuj84sEgRiZPFihCVp9whEpyDS
ZmjEiBAa2W642dEdDQCliActDlWe4sVMSF50qLcsTWeom9Q+8VbrlwjD5wLYDHOn
+OHeaYQJbZQYYl63dBHkqMLgx9QyUPXk7fkjthbK0bu4EXiBArtzGZHaUHwUAtvq
uKvQWda8LXazfv2yHu2vi/jes1P1/Kwr7TgSbBpUad1G4ts/7xdStJGR6gFWUkeQ
skbynPE24a1TlEzTPwMkbcuOCAm+UTwseE//bHLG04NvRXWDx1dkPWbynaUKwe3C
IMJdjaCXQ2SWLD+tPhslty3Pt/dIDhYHbwp1Mo5Mzk4HmfP2O9bpxjrlsbc9A85B
DzNS+l3HyCjPgwseq6oyFX0q7bj53WXrEC6rx00v5SYoGAeYwfY/7pvEX05ZFlQA
f5ORo64SK9UcIHTQ5UpnPvCecjvtplm3Jz4NeZ70WUZiWJ1YbCfrvbzwTI3pAqhJ
iP1EEi2JDKfHH9DOxAGYWssAf1eQvmgdZKSLVZzeDTRr8Quu6ozk320fvSbgedMm
d7lFmud2HpHwgC6JTUDWp1daZUTYB1SIEtLtuMjc0a6mj+bkTrLqLKy3NUQGfcrF
EGXLTDssFGBRsO7taPYMkVTAstPCQAbiHzsO8huodLH/8VEgi6w01NoF9+/bmssi
NADVnRYS9wfydNjIOGSJLCAPRcBWbyWn6berSz72tZFIS3wwO9B+ytH1NxJkw7we
njMgfSFTtzQyiCbMsTlA+FG5IuZzD/CNVCvXUYz6ab/jlb1E6Nre/A9ru61FUVKi
gB3PzNcvnVP6ArJLuFSj4DWyk/uavcSvUoZTxM9cPAGp5jasiHJIOy/MCQ4qTzo6
nBk6es32bxG/NSouh/x4stehakbKT4OdCFs2+18m27pcLCsf3/8tk9C+tf1uc4Rz
jvNb/EKjgd5L9E6t/bUVax/sy9c4SsSCEG8ROH1GMrJxl6tYC/Bd/uQGoY9ndWqC
Q6/mcIEVEBNiPVifTD6TNrQpk7v1DnbeupnQAQzslF8Y685C5uvCTiBPHu5CotL/
3F7WB3U2U+vZsioORzQwaHQP8WSV3zeuMnlTdmQSEpgAfYD7VrcEhFeUcHGvMPrY
feCNrMzNgOdaJ/i1u5IXHYR7TeY0ynv/wLPErBbQ7BJwp6xperE4cy2k9BALZKnU
20EAN+4URhbKJW0tF4dnbIzyMDN11Rv5FnONh0PBjh0bCy9jCRipInXR0uzI4X4X
AHZ3fY8l+hPbFo66KU0MUQW8YCO6tFRfWIF0rA+TDAjA2D8cTcalsCDtXz1kaer1
2CKOrBW7rhKvWlSuYv/Y4Rb5/UZRnNcP3Olr+4DDMGfbvyUKlU6Yglm6pqt18t7r
YyyKoxKfdrdYVaXUkPNLL0/Nq4CR1bu/CuPo9VI/XWNLuv9bASyaKsgdqO4BKVwM
rVtaVNKpC6fwDMJDzsYAJ2ujnu+GEVbOZMTG61QynVUkBLOMa1ErqYEWLapTqFph
kh/f91Y59S1+IRXXVGlMwAT1EMNa/nxYRTdtjxYIFnarlS96tYOQTF0vK69lm/pF
GKPE1qpr/F9au5GqtsN0mwWSTCQYO3xIa/jPnwaj50UKfcO0elsmmMSJdFngLj0P
So/iBRxY+lFrmAtUBN3MfXNuYGXGBTMICNZf9T5ivqjheExFmtVXP8vcEEy4Jqas
cUzawzJHQLNQtrAID7T8lsfa4Ih2ipUjH14lHwFjth+2kbuu/bmgZXiomGrYLEr8
Z227l/PzmW0vVbB+voX7hH1yNZxj1O2xT7HB7PkeCuhOPyGBJKqsiloYbUmQniM0
q14YRVjI4Tw5XsBCqlgDbXbrkHeU6tuchp+4aVkq3Ld7sD6ZV+d23iT/Nu7XzEIT
nI6Yx4kfqCIlkY2rj0204kguaScStYGDo5sH/o8w8Ya3Y7QLLw8wLrAYwimtpoIu
7MpDSg+qmTUKiw82KMfRPiJDFAgY5EWkMrqbniXSm/VQpl2HQunR7l1DX4KK6QKM
tNRw28kxed+ocFAmOhLxHBNF12SVoiAgc2c1shDf658ntikn64YBUeFsdIiBxYs1
sLUTlrAMZ3W4OWqyRxAWIHmfxbYIWRec5b6lf470wXrMld3GQ9IfGhE5AJtA679D
+cdXRsdZUiLt+52LcBKRJI9CS21MHoMxGWwS33154B9zFT1UyQEhfXZIOhddjNYJ
pgc/CugOXI8v6d2Ma8aMwXm/T+Qsm8WWtAIRygwZ69h5pXWhRf2JRI+36CQHWXws
2cB/swiDSTgq064oLDXWaWqNgUJAmPKv2ziEx+Ijg3iXDuvKO9sDC6Lti3mUFwZc
LbLzCOxW2QKVo+RGoU3WgscSpcqdwU3jPO/EOq6SlBV1yxl/4XDmCZVl/B+5tf4i
2CY+DBEAfzLYhntDAdq87uhMbYuR3cioCk6/xKKSOu482XhzybEmhdtpGjw0OnVn
2L+ETZxyTPB1aziNXxGubk99TLMKv5GfLEx9yTbRw0bidxgyf8YSo9InXS/9Gbbp
d8ApIolrhTkS13SJu319lEMCaN44WLEcRZIJyIb4TcCSZGF0JXfdh98JZumgInl/
0i2y/2xbe/+OnK21Q2xra4vfpcOiHHQ6HJmn8rGyY7RnteI48HAaeO7l/mj6oTnK
nIqs62QWiBz++aiJomnQaNMijFTtPi/Pd4VH0LWQpQlNtfDOVQzSpQAehJPk3Tn9
5b7qJkOKzgaIdVvEkgj4uJP/6LCVGPTx4DZr0DteRsPSbYgSH3tysUEQVBFFxe54
V8IyLMKSLsmxucvR7ayDqFu9GMW4Auu+esqYB3iTVpZkGmRKLTgCLO7YfKLM9RNT
y4MbC2GkUrfpxcpH8F/2hvu2hgby/ftYn92Fu+AxcIxFPQWSI/CtQxJNqOwnOLIi
4clkrgf3x40vhI1Ae5rPKrGKrCk1tDe3inpnECqefbTT5BWhSNziAGIkBd2JBSuI
gFL89LduFllqi4ZU3mjTMh3EeeRrPUyPvTPeJ51jk5Y/f7+Yq2Uk6+Jb3HtompDs
SPI7Vhm8hEH6QFSDF4nm2RWP/y74YEpvvL5YEmzdRa9Gw1YdFItEVkY/ScXpz5b7
LKZeu3azgjesVKtr1Z+MgpsIt/Ji1LcBMwtvBYLZl325yA/ghtF5YasB9Qn58MyS
oN8pJ11uICKFsFls5aSBHWgCxedoQXDCl2mFIlBjaGmI/rFBdbLoJh+qLYwrOBW9
HcpSpm6IEHVTqjWKR4w3SZ6zaqGqJSX2npHAAbwnX8h54rIUqU5f6bENiBmawbmT
2yvpz+y0Z9csVD1y2zHhZH8M7jU35uJTRq+SFXipBWHf8RPSOE9ZcR9P5HPXSJPS
WJuYqAMtipJhbq+aOxSKLf7vSkONidu+VF7EaDkpHrG/EBVARLpD1sIJoXg3VZP5
BOLkL8HWmGUDXPG7i38e/egLFurNcJIbhdZ1pRF5Qs72agqxfUfxfmbouPHG3qxi
mkNJ5bAte211BNpVJEEs+XzOWYVAUOxWVQmYCVnamzqmeMRAXPtTSikwoV6BFhjA
x3E4W0oU+f1fjINeTf1KCkWIVRvLKfV0/aXohYB9dlAmttqmsLRFD9I+cynCaBo5
RKv9/nU0eq6PHzpE1l/WKvylfWNJWkdEmpYJJ3i88LAa0tdqfZJqRBoQNE+ZYpwO
wFIKCFsTHUzRQCVchej9bhFR2TM/WX27I9InsMQcz5bjK0kXkAUI0J2dTXsKUr2b
6tvhNm1MYLdPWE/6DSrXybJraH1tbbzLAICAYgVvPc232TJ4BJvmGRYbKoX/qwRc
8pydIf4TncWD3C/4ZA4DB6EqgfBz1OGEYCaDglPkrhS1BQfI1Vl3rRqaw9q4koME
EC1qiLL5a5I+Bpe9DVwXTRtR/lL/sDw84T/V4D7QxLU7wh8CwPfdxrN3AL3Qq1Dr
SBmPjnusDTalkIOCry/vRhbjVQt0iRzcIx6jSsm/9g7tmnCCMbIXBE/kUgVpTF/r
E4Bhd+VAYiUg1Yhjj78SS5WmePe2C2l9qdTiUEXP49zopXwn+JVPUZL+0+NG/HBc
21GNOfnR47xQrLfLNlmHzJQlMu231ua3oHPDPmISWRZnI3Hvwf8hN5gRpT/wnYe4
cfNjhFhDZwxHraqvmpiTYn2iZbGe7OaPlI7/LOAcJUVBALsSSP59m+Cmq6j7S87H
BcEV/TavIqRQI4A+kca99KHz7zIe0E1wpnLpVRUdH1PGEnqf9AM/K2DTycGJtv0p
e5Y20UwNMe00/6HRXKrJxA69G4/NDWBByuRqUhGDxNw0YT/462WpPbtdMPPBn4jm
dBNXjjubDuQIifhb64NYwmgTj097GG3jYEPujx+vpxW7S1viq3To1g9pSJ0FFFtr
UlAXlhCvgESKijnfgbU/beKzfG3LJHH7x5x+NA5DsS0KGAvctH+Ippds31lxPppV
NyWjjCdFBevtCNwR2tc5nRJSspe/i4UkSUmHE9O3wJFgk106cs+XqMm3THIIsF/o
4XrhlIDErLN8IqwlQVqX/Cd/NnWJB484Jb143c7nlgkrmLEg4A8lk5tyEiOtmtzi
QGae/fGwtFpLpGw5bo+NJQpsP4GOwtLnIUiaz3UVnAnFzvbl+UAUAD4LcGvRR6eb
qNBpYvGJSu3yrIZQCOtcwhPIhj5BpRNWQgnjh+iof5sqr0iuvWRewPd6zQaE8u6B
RWyN4QD44TfUd0D97+qOM42bJkc6+ndSUURbn6n0vGvVDiEAGPBtbrjfKa+zBz3a
BQAhGyrR9d69Rn0YMEUHqbaHzm8qCRdBOr/lHuwVKt4birrGxu8cXToHutzOshk2
EgyaBspvyZ1Z3YdwiB+Y8B2nK23gD15KbF8Dj4dIU1T5jlBx9oeSg/rxnto7JNS9
NM8zAes+GClrAbmsF6D/XvtBEMgM1B968LOMLLrqg3pohxYelPqVKKDx0RfXGqyG
6XxIuxvHzc06UHU7+g6TBA6/S3TyQKvNbV4rCkdlX7wMXphOYLR0uHJDntQTxI3W
G/wUilQuxC+ntUwTL3BsnIs+Vqp+kpbrXoXMynyRCaARJdUyvN95PYT2GTZdCyG4
nuqTLCqNRIVCse4WUiOwvc6sLRpKUoY3t6xb/1ndIQQclKbJMPsX61u32parJSJZ
LnWy1/MDv73ONP+ZVgx2I4kAbavH/PL9LXloISSP7GtROAfXtmydDsJCcBti6nAw
+a4SYLXc10Gzimg7zsd2pQ5gONihptljiRH60221zsjU7w3Nwq5nYjIzfltmTQCE
f+SpUbiKer7eZj6lpLxR62flhV28qyZg7FJv2AX39I+tOLm0r80myDOcCbWp9nxU
ZjBNzjBfna2tPie4wOtFwfqvfPsBVjzgRx5ziaICDdabaM7leKw4GvCC4+wlz/zX
vVqRRHOvbTIQgHaCTpbJgvS3M6mzLTAH+XlgGmPEfbgAEcMQWsFQM1t5wVCTOXPR
hbV2yaSAckTQkvfOKrUI3HzzLzXQIGR4hTdZX9CJ9IPpNKF8DDClRBoVgTJy7Sl7
ogAG4y/NiyXHA4db52poFYw8QATtmvWeAuvFVrVmt5oD309GplaYtNCZekPJRJu1
et5rLJUlWQdMUP+NjB3TiNbj3hWju/ZBss+V2eJNgk3ZYrJE//7rENFeAEFxdFpz
CC5ICxqiewB6Tih8jGOp6kbbj0k45t1zpS6RbdVHwj0zgHAx6svM/UqVfbwf8X5e
Eie4cS1kPA8dZ72KXGRTj4u1rCQCNPBgVaper2IqAWnFZv8G6CC8yDzyvpmpM51J
nHVcdtms320NAgihQUEbLfURKSQV8pYTn4TqGSXJUHdaPoITN8KxNB2oQPujr/Me
RU0gm3KlQe4mHGdn1HNJLdY03UOmVLU9qY46oiRObMD+VqlVIyrwr0SIrJcggbnG
kLQceq00yMEBLlg6dulz/bH9yUFsyiJeIplh9mE0U7JyxZkZ12OeedeSlOCYeTjm
Q5UvZzYVj120vksqIT7YnIICWZnBNBD3OcfoOGEdkFlbX08mpTi/DnUwyaJ0flMg
KRSi5FRuQZmKE2zlNenjbPoWBnkjn0nRUxz12nSYk9V7K+sLuArYYIZ292Mni5H+
CjY2nPSoeQBgyyS1IZUhp15VmjTUxhEr8XX4BQ/4E7h17I+NGix0UP9UPbRYf23x
ob2aAvZZq/sjnGAKtsKNeAINiFWolPirYaHSeZ72LHrzXMltju6djE3BlitSChy3
+9LmlmL655wsAoUlC4aNPMxQNA0At0aN9rwWj+96PrFZKuFScf/iF+Mkw2BF74jm
rW3oUeEoKCZZcF3hLEAXFOYCg7awqSpdjIprnbhkHoklUtIKwH0vk5mTJBkkBHnq
V6VRrvF8M49cr2ESsxZ7MoEtX2g9PKPQ8kcgb+Sz92H7QVkdbTRS4NP8eA4qsbyg
BLAFo026G+5hTVMl0hPDM3N4V+V4ESq75W/M+lMNqfllTDPAGH72YeXPAsAeO3uO
j+KDysTcbrTcScS0Bqoq1x0KtOon+/7Hn6UqrgLcSPVT7iSxdWYGbrh9PARqUzCw
F/ChboAQ7k3U4akj9AHUHirwALSe7AxZg1nFaeMOT+N8xQcvva/9LxGYxWOJ+Q9S
rMgFRFUt8oVL7YcNXy/j88DC239itk0sYs2Hnb8qT7AxXqNyA6z3YtlsiX8DOl/j
nZCdFLl4hubDVe0+1EJmev3btbyp4XlCP4pA5DCZ6DSba8ruiI5DSSW7myMKPTlA
ucWFIdE4p+BpXty+x/QqWzupK6vUlwYhFQhGg9oiUetdF74bBOYOVPq4Tq/NvUGT
bVjuq0Va9FDiXim/YkSdyAUrpodOaWZ0vAr95R1lORL0g6C7kP9cWLKbdBSZ4cOA
zOI5OuzwkVo1lt6WB8Md5FhMX+x0rk5sLTazM97Upm7zi4aL27fI7xiTS8Mf2t9S
NwqxjT3xyB28vVcb1+zWrWxa8cA1zqrE9Vy2i+t5+neZmWwfr9tniWki6KGXXBrx
LfZwMckX6Z2ZQhs0JMlvXf5izci9QmN6qfPVgNzdyNl7ALMxwrW8BvIatp8cnx5g
wv22f4Gpx9HxTXZJ8xPdlgVDYIXWWFyxKUKwvy+OTR7YJE/LeeMLpWOThJHAo2hp
1q+Zs9zYy6s3KKnSINGgGMh4eQoLp+npjziujsA/bjZDQ6MBmcAKRrrxJKNM1h3F
82AOKTvlnS0iM3SH2RxLq2gReqbxlOePAJFDcQm1metJtj2QSzDJx4unr8Rmgo7y
TE7hMiebfBvl6xmeSwhIvKvJ0+BizXuKIozIqAuffRiQqyiA1cY2H6IpBAfX2kzP
DVk6p877bHvVfOi7DEZbNszg3Tf5Jb433IY/XHGLq9jJVSVJyE/bPYXu501ADSbg
MqUzPhdruO/pdiPl6ZYPBB9/ujD1c8AuASj1U0AyDnlKAdwkmrBzXT0FfT3AeVS9
JmkVFOk7pjXnCKUwTQflP0sCRsm6I/oFm0y98Ok8VYsj/s0lrrnP1FtlzHo7qG2Q
xHtCsnboXydYpfW/jUMiMY9FTcbvCAQDJPJnAeHamymHdMtBAm12ToczWaYgzXbz
tLMwt0pLuKOcTa0WVRgoHV8k59hAS1FdGCOKjyseLe/GSpR2aY3u0nv1Aw7oJ/WM
bhKNvbnJpblQsNhRzSLOjaCEqI2nGY5fiPes7x9ARjNG525UgqAigro6C23ktqm6
dZkRNQW2CDlnBrHtC1QI1GJoD8Mz6G1UEQUUZ/kkPeb1xFOafqOPYm5uldV+BXJZ
j4ThjfTkWMHuDDtsSVoJ3ASXp7asEfBX1uAkQM7ZNtQlFoiwX8VADazZopvAgcJF
7W1RmjIu0+JbXf5JZrX60aYAfvMyQnYlmJH3F5Yhe10uo15YcQiuBVGbTS5rgHP/
BULKWJ9VZQClC9od8JaiUaAmFVoCNenYtn+/YL1outC0arHyqQjf/s6zl4yDyaie
KmVMdcrO00nky2nfSkR+HH9NrMbM1cnQk/W96B67eE9ndwiY841bGy9oxYUyVUQh
Axhg9OgdCpkyJYJUtJ9d/SCWVpLQ0K9pX633Hn5mlVQUOkngNZZZzFWAMxnpD5UU
J2tOCHlcu0uytrrkxZt95hJ4G0RkxOXL03mzQt9/CPX9IKLtsLh+YP0BfN4wIYp4
NUxgGQdZ2+Td9JZvFKebqJl2SrAEKwYHaWoWUbe0tBLontVMi4d7QcdTdDl9THXU
Qef78GEcuuyABlAC70iWMqJWmWusbiL+ZiymoFuNXwE9Db3+wrEJqduZ+LX5iS3G
E0ksJUrc9VsKdQ55+02ttiAppj26x9GZLtlkYX37RVGmAiyWt0KZIoUPDHbzbIAX
WvSOjozcn0WTbOYAy9E9c4T1ylhIsPk0ybvfnTsB0WWvNa52ULZOgqbQa/k5tzED
e/VkErnNGwGH/12Zqt/zIELL3z6YOvfRoUTnEXWcki4++IjGwnfHFeUlmnV0XNlw
Lmoq/sfi58wdnvylFcXN33yQKQMJs9rkKyVUtoTsqAU08YDIxEl9xYaX8qkrQIXb
q7TqhSTvmA0vVck4Q1WH0eA+6lqsoKLGSkNkiEEURBl11aXk4KziMRJSs2qXJ1o3
fLniQ1banyg4LRUX85i/V4O1Q2YHZQ7dvMl0ZdtxX6wLu2hf5ABEHTwi0EqhOUrU
OWEr7aorGnZKx7L/QzajrsphkeDp28r6rw1+DU2zcqrl8EOOi+jX6HCWOodD3YrK
R0umYoI83vdaEYqgR375GYjDwLo1cRUMvnl3ar9SqgjXWdAkVFjMomnOU6CjJWH0
hVfeqymHF4HKW192iloFlACLt5InjJoYNcfOFvqB5pZSzUl04T4p0XgCBFneWvhf
PxicH1KoBbY57P2CpF4ZUOUWQx4RA0XaD5ndST3gjJ2FHp/FLkNPh3cNbAlixf4g
W3uB7AfUAoksIazwPHMo1BQDDINGKT0VxDSrdYot6f9W+ud2T4pkqVznKeFR2wqe
sI2y+6Jk04kFj+YmdXjRvspUtnPtI2VKcH5aJMWb5q0wrqUtQBBWNWnZBpuqaRjd
vSO3f/FoO8IrSoAV4XegPTGvW8/dPsDLBj7ooLthN4ukwn/Qj6jTiRaI9tfOaINs
ooiEBKkysgdwuj659DiTQRnXVRjTB+2l0v9yDa9VbtcQZrK9dvtKq4oRvmaAPFQY
vAAOlSdj53Giw4xu0Jl3fIr8kb3u36HIESltZyoGG9UpvfOa3LjrT9QbbdZAmvwD
XKnVuTZj3/qfPwzfz7Ue4TkLXb3jEaA9F9+nA8YhplTLuJYhgzCxTKaRjo4+VeOv
+zCctIde4STHLwFdtn7BeBrHoVrWQMp8TagUUVaiMWeaBW+mdGIYT06mLzhCb2d0
aVVd1OBTo51qi6Q0F7vwKGvQs/O2e5aU0rMXsDElfysZ4sl9bJ51PfCh2OcgWu+X
bDWw3cWH+79tqIwVY7yJqpwi25pjp3GqOmhNrFOpxWt7oD1EuGIMdQAE11mwwPlu
x2QbV3xUDcKhBfhGZMCtS6th96y2UzMV+1rnibVtlmuOCxWhWh1hzfl0y3OEaBEU
p5F6l4810pL8CtsY6CofLgef/Q5XCxLNO458gr/sX4hV4Gqzpxx0IzQ/c6aWvzjA
unPQ2/DCrPizknBhyImvI7ObPd4pqJtDthR376/CANZ4wochKd8V4K5GXdsNQW7F
jVczYVC1ZKM/ZZjn2CTmjggHwYku6hIYw+ouWB1ED+UkGybVXVM1Xui7OKxc9yml
uefdpJBS0yh7+gI6Onfg3hJ2w/8b2n2rYn7sZSNVu2l+u9x2SlBM5iVGzE+tP7MT
ML7oh39hzgv613Y7aFb8sdZtLfJKNtapp5F6OSmsG30+vECxQUrfM+8IpC+9TzPi
02cWm3QhD9DF1x+aybEkDi4oV1eNJ8epbbDFe3WcdXurnZcwp2STCPNlPd8jxpcw
kV4jkJO/6XX3ApxmPhSkS9DT8fRU2oM1Q9oE8lApy5pV6gpUtpFmiQZMifZ7y+3L
cJRJ+god+UJTw2a+jYyCNfbBCbJe9qxPieUTLERqK9xKNcFdkjfNYFY3HqDqY5Jh
nKSluy+Ntkflq7z87AkLenZkyt+GIXOJjfC+C1mTHx4Fiw6ERLqt+gT4gionniUT
WaOfYn9wrFkKmsfbWCzkWox0BBOX1oEJGTFrO09dkuh/lh69RaNW2+cRlFY98Bu4
3QDDQFMNG5h8FCP6cU+C335sWxGBeJvharSJIRYu1Lvxly2emb3ezkzg7xKGdojH
DEareKxHWNShLEwSmg16hIN5iJxdfR/k2LixhQU8h1flcgFj2Q81jpFDN8WylKFC
+SjOOeQXZuE9BL2iKPp1waOPOAuRV0CK4o6HCa6wZhEINREZH8SsulUSbvB4djGP
dS5pDQJB25P52cHvw4sUebCvZ1F5bYC5l2tsx/00/OuSrnd6IptzJYa00dJYzB2L
kjBx6b7aSWLMs1a+ZMYTve+BrpXMIelRHTKvhLHeXytX1sKfc5wAeg0rCV6R9fTv
rh6N/GQG5ZKZLQW6YZob9eYMZHykggVgkW3e2YFsPcPO1XLODz0Ag5UPYOMMoSoO
U1HdlXsExZE21LSnjVpecLYnNCIAZkDnReJoJJcUpYnv9J9MBrw1dzVjL2Kvu+3A
hUHlXBK2a/Qlz0/6jYWZrHVMxU+WzUTMwxxAnmDDrkYDNvKKneIbye+JSpD7ajgI
3MWh8m52NK0rRs4/5zRbPXzfv4HpIxZ/hPWkVnPuxMetFbe51JS8EOPPWb21w85I
Y59H1SrTWSrk4OyuayD8hR3i1ztQh5EeC7pUkGlAXHaSyMQHBc1WYmg/VHlhpAVU
56pdsTu9YLSiUa+eQUhKG3oXkmUbxBMAGytZksmQo30EKHjD0uAvZ/whyrtHqRqJ
98ct2E3pZKiPQWa8KyH/80KGF1rBu2bilBleIKk3ioeXgNm7m998FxeVEMdYXQrz
MaTYcPOIzMPv5ZgDKAZdzzS0wunMWlWSPBtBOPJc4YgCf9W6PgesX9i/Hcjpx1oP
8GFxOLLidz2OPbfknbs89VJNhcfaGb9WZHNNGcC8Newzr+WkpK7w2goqfsdgezk6
9UwGnpETdnj3niPbl9B2fmrK7hDxxQYQdKJxbI77zK7DBduPU7fXHuYR0hj4LxhO
WiDZjEE4U0P6ZWDFREfI+ZZlkmk/iD/YV7GaJr7kFDRshiOFWX7/7iK6SckC3PoX
ZGmvxEUPoKVaksIb40uTwS1CwnJ45YQt1HEBGngnjYFl7w+rNynEnHDrutJKEpEi
JeHCvbTlyBbwNzYJJJmcdObqJlF1x/loRDGuUHV3C4kDC7y7vAtgt+6sfp253QZp
eOEpkyaTD9qE3PEjmywQpSWeo+d88ScDXMozkOR3zvgrr4V9rG2j29vNmZuWSFUP
alkp/xmp4EXFcC+zaFsAuNS22E7nkfZkzsX5GxlaxRs+0RkpAO+IQyaiFA+3RtQW
8jqeoPYAEwC2qSwLCTb+mtC0G3pBztVSYvvf0UqEIZ4rrqR5xPQgnPeo4SYlStWD
J55KJmH7B2AGQko+wZmUZ4gm9zp/Q3TqNVYt0RExT7fWSjEFfKBITA4U2Qsgx4to
p9c+sqggG48ZdtkEMFSQTZj3jzW2es4hdcOPUCXhcEK3/Bs/FBxT/3crX4sRmJW+
iII7T/h24cRJxFR+kVtS9fSrsl1S13Oj2hg9uY0Aw9gTA4aZOksX17mtEbUpGRyP
W4JJv5cnia15f320++MabItTCRIu9qJCqyeLJg3aB6/H6tki4jJkFTnFfKttCxIK
s7aPvnUwjkNGzQ9+VUxe60ViVAAmVk30D2+AlsbQna97G3/blwqI+oi7ZRpeHFoM
DVEFw2xymd9qX8OuD/SvmEL2/go8tIensVZgJhS4TqV6w2AvoJpsZGp9db1PEEB9
4ceRFuyyNEGqoH0ZrhftlgZuFUzbz3vR80m6Zwc84uletHPizxWvhzoeW6CidhwT
ldP9Pv87wNIqZ3EOas03hzIBy3Sq0shK3E+j8jy3gc3EaurNGfK8t7+voLClMupU
ZT/pl37Q7EkV/hMXZzGssWg4daUlqx36jC7cRQQYTJQBPzJocSgkcmdvYpFk9mMk
s/J0N0Svxu5xpHNswbozaU9i0EOzXXsEpxtjWqN0DcwRZzjmmiYUlWAPayJDfAWq
jW0iSGdveEVNadW5HiNNpDxjknhNv/5Q/BIKzgxgUPm15ZXszhaKm6aMjRdF9156
TbL+ImfPR7uxYKyYvjpz9DkssRp1EWcjogW9ROEep5dAqBhl21VK2zm5RMRgbXu0
jLbadEZ3ncz7yKVB/14E6xk80W4IlGGx9MeDm+1tl3KxnftwgPdfFw/fL+66LRxB
8AYORTclfQi3mrDYsyroF0q+7qFMmZT+UUpTB4ftPeqM792luzKF2nE8qhQBSTSX
kx6Fp8EIwW952Qhif+OBKzV2lYVyXY+mcJlaJiER/8iD5Lt2A+1zuWI0iKNifGxI
JGj8adGFDfQ51rXlXxTcf3KOEl4mXIJOOMRz9nsomDnlHi5jD1eE1/raLZ11LFhn
4Q73ad89e8gCZM2nSQDiRWMz1ztN5c9AnYqwDrGvgrSC5WUSdwaNhzrO2m6jdsxL
GRr14He6aHZi8EecyvRmHq/F37nOYku310/sb6+grhLIcd+Tpu7v3bg9qsvTmyb2
xP6M3XcIc/6SqpMZQkHKKY5IR4uyUQ/Q3628CjRM4VuM8So1+9RBEkIP6dRZmU3c
kWz0sFusre0InGj8/E0J9h/nZRLREFdY8T51J+RGr9PsWlErK9fCMkTrQnoxEJR6
E38f2fFBKzrLQ6F1z2Yg5r5vXnULB0XV7d3dcmNIHDv6OVHu/8sQiGRJFb/MCMWt
pVh1dbjl4oxdrCNJXK8/qqqmDzqEZKsRlWeICztHBrDkTKBw2c5HlYOVVSGvwDT8
Sn0IwgGDVDseUbhYyfLm3CrPc8O0v4TpxZSJyA8/XxSZHH9rUQkodB3UqzxwJYCH
kR0DQJ/mjmpDs7iVx+ckqcSA3mcsFRsTeaoDJXwY7/2IEnHnLFzmSIpEPe8+hclZ
lw8Srly3XHtfOYVZb4jpsSGDGrWwM5WOU8VR8qWaPIseHixR62+9t0lUY7yjTDny
mQ2l4x8oQpO9xAFOtMKmn1PR0cPDGCP7YW80g+OtUbFRqoiPJSdARQmPfzOT+XkR
cFhRYnASHKNrDa5gXmwo3Fz/b5I9+hiIcUB6dhzX2YG2UXWc5lByGvEu9AIhmysJ
EQdwYqNzIxYhJfkutcRwj00aaH7wRQEEprqxWP6r5DRW3DDi64yP9nUjLlWo7tkR
mEYzcy+4fUZnyciSBxXuAyjSlN2kdiROBRmOSTRfrKOHVUVtmSWImv4Lf0yEU/2a
WKQ0Souc7FcmuMy3MX0IuxyAryv+6Vy0TPQgmQbCw3yqI2QePFw8eDIWWkMlldA+
uJGBLaQ9grJ00z5RBYvmUq9Q3Flsp4IpfDirpOIAIwhrBMfJLCUWLVFxYfcIfaOa
7WYud1eNsJHkpqnbJbujX+b9N/tId4ZUfjcMGDljWhIHU/PFaQJmBROLJq21x/DN
bZ1ej/xMO7dx1jnYn482SEeLs4SjyBshvHEf044fCbiI4Fsj0F8w7bEqVo5chkHt
EEQ8mNavi+OOxdGSxcIuyht81EiJuS227XDjHt/vyOhtnkwL9PBCDP/d5nxxhOYK
/bBWFoMG8uEtYYMFymAY7oetPKDrI6M1SPcSRnOrxI/tSXvzHpBn35hus+PUicvE
iaG5rB/LpyV5eM4Zdva81qT3+e7w+Zmwisu6l8u/2UQ/JITuYDQ9gLegtsxXc3KZ
b/o7Pi3SpyQA2FmrNM4LeV3190kgxO0JDDEWGQYEYQLEUGUdRi6nMpvN4p9kM8PC
LrwPYX0/lQ6i7PJj5ZT+BtkOcB8agW4RBrK0YGpyygjMA8n1yITVDsIaliDMCd1j
1oEjCWLLth0JP86BmJw9/EqhBIYD6r1/SVZjrYj4vIsGg1UH7NWAnVf3qr4GYAyx
Vl3H507p0T5c6Zz77O9vewoox+sGT3eatL9ALdUWqTY/TmVWi9LrNaQSK2GiziLe
/hvXgbd8Olg7BQaqmXYcg4KOkalHCZ7uHupbuzHpUfwdjrleXwkbxa+0QCluqY6k
qiupPuPnrSKF1LaVzwN5X1eM+U61xzGcefo6auEqqv6GNUr2KKkwyKEU1qVB0VF2
s/WMYvTBH3Pg1mIcN8DWvyZ2C2myCy5XFa7BltiTHYo0MJg8aD+03g0DbGMGk3AE
g1UKAjZ4PrRmJGVyL+fDUunK3dXTAspIblfbppO3ZmjI74jKstQhJ07wAvx8Mpgi
AEKBLUYuIy9wkcWW/KK2v1MQ3g1DfxnPMtB+Qo3QpPL3/tQu7d3VJ2Bk0cdDNaI2
BBDhMrxLvcSBFVwxJ2Gr9Xsxhg1Jc4q24nERko9khFt6aDwZ9Nv6cMqW5IjrTJIy
wyxBFEeu/M8V4FSJojNCi35Z9PwlrVtDm9B1wkI+U8gssvID6sENAnhVEvaHGRoV
6TSK72gJRNIyHNHz1C6lnUYIvvwW+/lufTBOHhhTI5RIcK9giEXYmLo3eet+KhNw
XtB3gh8wjUX2D9rd1dldnbLkux7Qiyk6Az+Fn5XOwoGplPMZNPBvKari2lvQ0PFU
MbWbfv/bpoc3MJhrj8V+NWNbq5S0mw3GsMcIFSjYhh+WmmlTbOKo1HZTPX4MArRi
xAge0qrU3NNyU5YyHrFt6jPnAqSQso1VvjNdJAwyWaY0/3Qe3WoZEYKH6aqsVtvm
DmcTIpBOxKTZs+m3/Fe2ysPLowmPKbt68wWAsKfuy6WDlnDESKy695UJB3KLcp2y
/gXrY2FAUq2PF8h/9Nm2LqCs2z1ZWGxeAL58kyEAQjelLqM2eOqGvRLKAmn2ftAj
IPFORMcSvBP8ySOjLI/DiYB9343SS1jiqwwX+7/A11+hi03JHtivxe+oQ7g+QSOT
Ln13J3ShTQmvZoEtVwvJ2ryNbw4rsRLLLOKBrfVZrXjQy2BoIYFH55UZQBKPDV/b
bLlBgK44V9l0K7broRb0H4iJMpZAeXy/Y11AbHwOGPUKKbkv+sdRVjgDLWLoVtf4
4F8gAe2sScEWxmU9q48HZSAgTy5cVagcbVHRM0vMx7ZqIpcx677jhvjDBQ0D2d+R
fwv1gfLIc4DKXgPMNrJ0UJdfYYezHgLt05huPJIcvg3WXxZcbn4yEDZqLCAjfT/O
0LZ6v2P6CNbhmlSWPo0gOUedxB4yBHYyWGsXl58A6zTxjiccsLSjDjvmmJFitlNU
Y0rVoL+3qalKlZ22D27HhSpW9zVFdOyyyV9QdtmHPMf0FClCBZ/uHrXi2wqr2jKH
Bmwa6NIBwFIu/w8lST7ES4o7BBtHFY8kgOK2l5HiICHJpHWE7y0jFdgyiphStXYz
ou1IFX4ZOwEeTf4KmAdfyCK6MHhfp5mIgB2d7hu5QGkDL29jdhfGC/WQLxJ3zUzc
jLBANgjlwgdiQPVis00u5p6LUkc+v/CCkVjcPhbBDtNPYjurVMOplFDPoCdGlONH
xNC2iAnPOq+D7GsyjU4K19Ju+xc4+nQYAZBn8VmJ+GnrMQuTFTLkCXOkgaANbOwJ
/wabn7q3XWZ3nmVNOBhoQeBk7ImnpIlzJe7wB8J5s0TkxVHQ3J/cxAr/QRBzH0Fo
fs1rU+Mzb4RBsyT+C694nxntwDD/pdaMlj8EnKf2frW5Uf87yq5KFPAFd09XpPmM
/rFfbss42UTUTd45rpoZniMF9HjDfBaQkkgzsyelKpAlhPHBQK7MU7y70+91JKgo
Qza05xNpUuwQETxRRFY2oI8YW/5QOu+btrXW0sjjaAreGgr2oPU/puUtg4UtJSx5
7rjISuvFmWxsFBlij+qeFTJnkrPAPuz/oY+lM8tDOdn3wiAmWZ3ssUZ2ZPbM/jtT
usw4N4TZdm2UoEkZVLHwtOTh/YkW4AILMPJeg3LeTMarSpykFHk57JoAJXs6p1Dc
WsF4R9wLf8teNIFNODGXKbwrS0lSYaEpK5rWL1QnN8dZCJhdU37oIVOkjsZ2t2eQ
CEXr4sN3tzjeOHZqQsUW0s91LP4FTVKeokNJV0H4PYyQYeDsoDH+m2ZqofaKgVqC
IAVNdxjwgcSxhr9UZzKNMuhDDz0wkqYyWCQsal+aC6f/lqXmCE/gasEVlCH5jUto
4Jn4OCpXrz4WhSYTzwv1xAKjNt42k7kHZe6KCLBffvDQ8zIfRzfUnlAGHjOQ6e8e
OBHYGdibzopTB7q7J/TozsA0bl0x5RgSQM/L7vnCY84IMQgVS/nzwPY/GVIB6+WM
wn/kY8kJnl8cG9zKyAQqe4LYIci8eSvxKWiB3D8NTKp+hFt8+jECgFNPbDqAs9s6
JYIvZH5yRwGx2cps7rFLUnUamFmX2htsBtThyimg4wc6Kh53blSexePdl4362bV9
R9V0D3FxvaRqEa/DS1AeX5idO4RBedRaQUGOAlt1SpiIYr0cebBwp3nPcSFnEITt
gO6Jt9QKg3bDLfbSG+UE2xH4s+G/KuJZnExtrKfrRAMYVxTkDqHjcWQA3Gffd81S
beAMQiMdOTM+gbvInLJHjUbOUeHQhLXcwmZh532VfsVDWqF5awAM2jLjPkbrRFm+
sqVZCr4f3o6qBh8wb4qHxSpoiffp74z6pl/R8PAxF7MhEKU9VPnsJkqD1Z5tojgx
JHFcO3aMYYDGxfmNDGc9RYjohDt8ICa6/y3IACU39IBtKkoPBJOS5IYK6u6v8wRt
34IWC023kTvpFNSTp7Gb5S+o6LqaS5o0oCP2NjBdLmrOHXx8FY+/P25OZ0GzqxU/
15YWnPbuQRyzXlPj1+4sLBXpJQAgC9WXt56BRWVZ7vyOJLsKY4avgX8OCY8TAw+k
QtebN3CLLlvjtGkpxYVxxwC3EkRnh1swamLjH6mIQ0jCVUXRIA2j+ip+pwVNQAPm
RZ+o8fY00iACIxr49Ot0H13EY1NrVLlbkbWfap12Zdfksyzn6f65CbmU4m+NZeMU
fy3grhDMQxd28PUKLwD5gEm2cPXCXQJzxjcQy7RzqO/cr2iszmZkoxWTblonl1ov
IYWDBEx+t+ugkcurVT6dngobTLeVLjDrwq3lME9ULeaHcBckwcTdV9SyoLpuOjsF
7UO84+z8xMTZwr08p+VKNKieNyJ05zMFRN3TLYozYruG293bHKJWv9Sal1+OkBcv
yVcW2/eAsBi7yEIYj9k7MnhtQZOjC69Hv1XAx2m1N8KUniPJ27hTM37OOGdPrMcT
tS/ubzNy+hncnpg0f4pxjFzxjLwR/1ABKtU688nJoNeBzpF7J8Drh08uE7ss9/Ud
PmG4CS7kwk9MP7+OKb1+bHchW2x3HqGD6/vJIto7bqDc/Q1jOjUT/2B5IfKqUWb6
w7CjBtg7cwhSZq3A8OIIBqDp7BgYrsfrPa9a3FrlbhkAUzeM0CiJD1CxNsTGloWk
2nh7KRLx1qHdZyLQDKCnFcRpZjaoU9HjPbVWuyM4nu4X9bI4QrnPYNOsJqoJVowg
C4eOkkiAxT7UIb0/wFVF4dtIXi6TjQcMUQpW3T7MpzqkNe2f8A0o5Nw5kNIZKAzr
T63lbyjcSfd8qpWOPZqMmdGnH8Zjmo9v0VswNMrx/wlD04E5+nqalfRePIwaM6G7
C2rIGMMv6Uu+VLHq04XNpWKr+qfxdshoSRGomX8QGOYzE0xINWaodN+WXYOPpYk+
wg4ZklmlbY4olOeZLTfJhTGhTZViSaiCOebBdwOlm4IC27OV3rbdvn/8dxnh3ant
4GwrSDUZ89ao3epSpdXrDqiz6/335ukx2pwJlxrK8KwRPBDJ6Bb/V3YSadKmnOJN
9OhpQeovwKw70v9pw2g2Kl1EPOHDGuwylJCbG1uU4Lz02hruJ5vd8Si4aNwB/+bN
JqQ1+aCSLZlMOhDNloeEIArBqvCtArLjN/ABpazUOOaJHRZgp7hTK8/SmR1pWyay
E9hJbzCYKU1uRvEGuac/Ho4oy/1lTanVexIHybSKH/ao0kruvvBTfceiKCVnWw05
JzLl4p/fQW6V+ZcIAGJX7OINjAFgbOOM3+hKGq4Rduo8JY0ARQOP30g+4W3sLOly
aJLZw+aIegT9yzPnebldm8nSWB3YEhyeyRYBsKczJgiqG8CbtM1a0nAGwwPF/t/3
6lTGmp+7R8Zm7qQklX+AHlpagkMB4zyIkeU8+Go4dIWD7sUVg7eHmZdD3bWw6jmL
HEPWQ0IXdRnG2POVYU3GarK/uUaYk15SCv0wNq51s0beCKld9UqAxGt15PlS0pgx
9LbpHF/CWT5cne/qYJhq8Txg/6F0jbCv0f5HhMWIVAblJhuqa06KKX6PZZBxUabj
xU0a4R0ibFGgSr+uJMqZf1K4CLpq5Np70cm/qdfvJ16UnIAVsiLFB7/JJzCVgQpk
uSuXY0vw3SbXuiKcdAXaKCsl+kYA3T1M9ghORw8pNWlVvGrF9eHyyfyEcjPt2yRv
TlXGOHNM7zv1+QHxmI6Ej+5oPQQyXRBHmOXkxrmbkDuozqyKAISEdDg5sPP+aqHb
skiEOciHKgb0xAc36165hqGjpYo64RHUnrCAbT+WICZ3NijxmFxz1ahQq8Cx3ZPS
LF3OKJPIl7ZGVA6GKD4aRruhxrPy9/0MkFEJ0WB0R7uXuFLvcI0DV0goCKq/fhMO
v/g/Brd6nfoYPoMU7zCTSjoFxYydTFzzo4xCAq/HhtqubMSmBqAw/As0PUzM5TYt
XS80ULszXzKaePfY053/D6AO8vNNIVkXyr+WL348wf7P9JHtkuC5WDr6GbJ/gBGj
HRu6ZjCrFPtI7lDbh4+r/2ISCDJVNllESflXnKCI1QXO2+UlG0ROKX67DSbXgtve
AV3waV455+9HFb3+5roaAa5XROkbLvJ3ekkT/WmvCAxSr5nOEQszYJzLkKU9WVn/
6TU+PqZRt79gYH5m6J1RJKxkRaxuoPOc/XyklKwQfiiVLCIpka1Pv4IN5HDcr3kL
7TfaaEHb2LuHs3nCQLww4Bq4zcO81mFzWD80wI9BJeGqPmr7qJMa7nlwvVgbG/CX
7Vd0u2m3A93JASm6f5LR9zR/d9Qz+wmF0+VaaNj48Xb3ZxlEiy7uHo3okprDNKrg
EvIzZ1A3NJfUUUqR51RycVyexYsAgiRAdLTpsdmXvASz5zwfpE/ZH6NYkF6ZALvd
IiLwjyLwfEKi8NLk5DKXAJqhHrbudizRvkE1RARlrOzpoF03+o94fGEZPx9Hf7i1
89qEDNu5gd8hqx2OLrlsQSA4ehisE7dtaFICmdmuLFpOXyIrr8vlM6vnoslMUfhO
78YEP+lQlMnzf60kbp+bxemmu46vpCiJcxRaDyxwQIp1D1OPpPINckLALDPH5XIg
jENLkZF5olOFIlnxJxUKa0p7cW/kGtRqSfImYNutmoJoC095DOnsgZTns/e9DhO9
PGITNIELu2tr1thdBUnk+uF47Bke4FW0Praunrt0NtI739LPbEvXDXLhrDGluhC1
zTGhpLN64hAXUx6iPmkiI7EgFU7FJlK14Dq343Y5V70E/jF+Simrsu1kW3C7hSOh
+WFBX5G3yeVy66cG43H6ZtMdB6UyXX10R7EXwH65LZXvqKSOeVRwMb7/vIEL4SZz
Cq7oYQNJK6/kM4pgJxF67cOQJuAqZWei4JjpUvsqE6bzqZCnn0e+YzthAsfLerQr
F7n+Nt5IhbPR+DOpFPEOcfo6IX2D7pdz3FF6pd2uucTXUQdVB6m0UE+0pCBjG09n
IxDD/681FJGvIkrMbh3pU45/6Zp98LWs1x9tuw6MNzpbYi0d19EWFaTFLZAkUyEH
oeEKdjTx3SYjmUUzMSehd9bUM7JpunRSQ1yt2jpZk3f9+3DKCZkihJqMENU07QaA
wNqDhA4w9yKmxttN4UJfNb6rxIYOI8aq+XYW738lU4x9lYFAJQDc/9+kZGYMCe7L
MVvnuWLohCvqzDSUC3xzrL4mNcHmyjxO5XsWaNGQmM5z0/k1X1q+cawK0P5jX4lw
rdSXL8WHkEi/UCCVx2yL0STG1A+oNS2iOMUQAzT+lPdt2jdKWxFQrHOJ3s1L+rAe
tYGMy9d5vQHHy7ckYXtrwkDJdAcbChUb3uN8bk8Y05ctmfuVP1VnGxRNcdR3a8p9
HFzthj4JqV57bfXG5DKLHcZjvpsOWSMPNOyLylZ+1nEMOOEyfhpE/+wi66rPjFOR
g7f8MV/4RMOyb2jpZyfXGCcYjSUWg3NdbBph5lv23oO4MLJSB93QDpCMRzpqN12K
E3HyXMwLxKUUEUxi+EBOJqCiJ2mW9gyHEc7+ocglGZyXthPT2RYEdoo5o/fDBtcV
l3Vk4Bvk1gpyfJSafvWrkkAEMfjQqAhqOE9SlTqj97FdedW2gbp3OQl5FYooQe1r
JBuzGAQjctbagGNGWLaQHTiyJO2QnM9h6ne750aX+oo37joyrSXQCbGAUi/AmdXd
HxOXGbZhq1KeiSEYFo8CqNIUIJWFtmlgsI9dh5iDcfngDb2koJnlGiFtmhsjGeqa
seCk7xNo4b9wBjGfYIxiCnKTgdfSj/jSx1+70pTlGesQw0qUd+klvcGON4y0MVhW
n3uEoAUIT1vdu12DguTTOoo+jG6DRJjG/IZsbLZ1IvJ6BHHjOLR0R5in/bkQvp3m
nhMLeg0ztqytdFC8xe+oO4hrmp7TLx/Md51t364stSxXab6j5RQqq2Xvb+54sc4f
PFi3WJ8mKF8rbTo1YvydCZuzIFCJAkRmLZuSow1OuyahXMFQHEakpS3Sthu83Rw5
z1ZLDvUUnEXiisB9dNKejejqdw9mZtA6h0kPv5NOs61xjTT11hcINwLvAOFaL8F3
42V/VYG9muoXZrRYkGuSGuBpsumzrMFTpYMNUQKnfeXwLXqBiUl0bNvokFVktIZ3
VN6wo/vnRocikz7VdRShikA/Ll7jovkfWu1lu0n/G/t5eh5inKqH+CemY1bp0HkR
LLg2XeeI684Ihzq3rY0j+uWzsX8IVh1+RFx2yZCa0KFHh//SQypby0g9DCs7GSC2
HqKEbN/wmkqN2m11wtfbdjMVnbWLuDhMQ2YKxRtgeNOZaU7+s21VbMWFYUuGtC0U
0SCiIeNrFv6Q7mPB9NdYXoh4iCnjes0w2eyVKs1X8DmKtxekpZjmcVsWJKVtldr7
Hjb6TeeZ6RS4mEVs6yiMOui40sKU5WY2DEVXfUs0pPfHxuB2g+KdLJMyaAT0dcXS
0V01EQUZ17XPdmWj/e4cJ0uh1fAbBMH+M1TP3vf0Wf8LFKVBv9prNMfgUFxR3leZ
UVMqPJGg/+7kHMXm9S0teh+NKyGstAjU2KuTEdvHscI3zTZUq77koUDg/XMcByvU
QL1sRAbYmj/dJ55yKxtEuDNLG45JDtdEDRkSCfiy4v9V4K3RMFio/LokNvePw/uu
ICQuM/HlArQ0G2gf3yNugXWu49NtFRNuyOCgdWn+menQfLC7JBzQogiEHQPUl6m6
b+zS5bgXTIta8qxpceWyUC26CHTNEbTr+niJplz2P5Qd7ToYooeN5xKHs+gxJZHz
sKojEcPH0NzV9wLnxn97+WPYbar6/SkvuWxqfOaT8qjQGoAMZ+rGxPl7UEj/VK7y
3J7ODl1Fe5vL954eCInLJdKter9nXsXSoBkYsvNKTy5ecf5TyUyKtwRkzhzmIdMS
jkrDwpXUIR0AoAyAIfb86Blo7eeacIm2CAXHidVyg6YiRfCOKVezFMO/34uCIEkg
Z8Z49ZYZm9la19Q3vGs46LMJz8bKlLqbEmB7o5CgkbQ1FpE0JAMFpA0+1xNcCRTE
Vx74ZbVYNc0RpjkKKCwb+cudWStCbSSL0hH+PlCm3ZLirJMMniaLpQ8PCBtcqRxI
6jcyeLcdGxqXcLIkO8WRsIZ3kHwJXRIGjqIaqEd7cyDMT3BcjPc98OFPmUDr9pyF
pD3q0FsKIb265sGoNN4gpQGBe5CAC5G/Wle1YYp4s8BSTBeSN2ThSL3DvcJpCOtk
XCcBWWZ7S718aUGhSB2qUDWHiQffO1xMLePzHGueWXTYiCVdfloDdHSJeChht6l6
oCxkZKI/4zkcLqfbG0iNX2K+mYxFZAykhZjrvIsvCJ3P5xsFqhoMKGjd5P2OJOnc
9coSjiB6vd0jZrfpna9ADr7D1JR6RuJGua50nqhT6gy/f/+tfOts+CYoZHgI3RcR
nbeG28RjzbTa5moVxrYkXgJ9ubLUlH1Iq12iybIBEKHppPsUXu+IFdJhs8dFJOgc
NW1Z2qhAOCvaAyRB6/77ULNFxBn8juxRB6Se0yEtppTBIRoYZagcwJH8WvXM3eLw
RNUfJeBDuycZTateZlzV0/n4Csk731/M7bsr3t1Bvj8m0bMzVfqZjfLfTFw5WcTv
co5mbsdjXvGX8OcQSYhBQjoM0c0/dr5RrCbN2KupPRtOA5rp7dvBMl6pNUSsjSF0
gqbda401O8IKVCkarBzwFZ02qitpnj3HzakFcCLGmulz4tJzwvx+EV17EGhWohow
Yl5XZY8BVAAQX7UmZbx7xmecWjhsa27ZFaa8WC2Vu1d///SonHx1cd4oKnuKQy7w
eIsIdyyDiY08Ylu3k8D8qhUQ9ZK46Aahfe1+bIPxP1bgoOBwI45BM+Nj7S4MvCEf
Y3ZAh0ukm77xI2H+xta0UWTgoJafsdT/h/6cTAqHVir8Uk3z4sZE36lzZxWyOPdq
Wo5OwkPoQCS0TRtdHXIWPCL6rql7HwCe8OAEfrI2kBi/JY/tk3/a7o1AY7sxLwqW
DzO01AxddFJnqlZCyDPl5/iWN9dzB49PU2HCTd0FAHOXnrYhlSP8dIft51tXkLVX
r9kBvtJrHj/ac5T1Afe+aqJOCCctPiXp9SmWye4tl2RG71IbT38iiZi9VHm239Bz
xtuluekAePIkD5ZYXb7tNMmkteLEguWWQg+r1bm/c2k+2SDWZ0DPHzwn+lYarscq
8cKgmq2uTU+zLPLsmbXcir1Youq73h3ltpy4sxgZfMJhgFw4Qag+10xosSL8owyy
YTxgVsPY8Nf0fT7HI8n+07ImeMRMD83MDyYpJvz3CHJ9JfuD9k3Axb158LFWLdm7
4k1KLaWlLwDFcvkJ8h80nPQtV8bN6THiroBcRsJC0CRY/EBAOB4cipDts2+09eru
1DfIJmYq25tpDGdzYHfolmhbn9OqPjy6SVCjBRODv//sDXsYxsb3+3KxFJrHeEcv
AgbUhWdTA8y08E7pVHgyMcj9wg8fYO8ffBZdcto7XVSvNudLv72YoLqKRkcMEhw5
1dVHjgPZqiV9S3h67k5tsvlI9cHaANuI/4lBFMY9MbcjJrhlqqOWE2D1/wkzVljL
KZlUQhMgBOUK0RwDWqKOSv9D8X3SFPKbhssNRF2gKF/4KP2LRE77L7/2HFY+f6Pt
7gZHGSMz0ocghxuB4aXXvc4tMrXUKZFD5dCZUS7fBy5SV54hdK2dHJESSliVY8Nj
b3RZ/jms5unB75Wt0siuwnoNRGhTCwcUjb+Tz6DETLCn2kG3m3WG74Q1qkek73by
1qv+/SatVScgZs0wtn2yFejdjExEZBKP/NIKowtTBhnXRxsrk5y3XEZcivmZv86q
fYPaEUbNfWUG4GBkUTgcAFmXEignWV5JOrCAzJNXCcslgtHgEn1bPpQwgtFKGSt1
bOnOX2veIEyWUQoPAdWefUANv5IGC25zBC4yxHjJEnoyUo0jH/IejycWpJmmKENf
GXie2LgVieGYnDujq275w8y01Fj1+Xz05wmB/Hm3Kb3/i+FM3CW+dOOZ5NTyPMtC
DuutaZBuEjIJZrrT+tjZi/apFCitvf2Jvy7kL6/AdyG2p8XqY04/uUtkABCy4j9N
OLYIyD+dFpnVeObelRv/hp6Uc03ecItgZKNzbZQVzS5in0QXHAqn6by6dt0+R/KX
Fu5pfLCKehWexrv67l1LA/gBLuH7EdmIBNw/dNF0SItmGDUpLnWq9QQZTcrWwlb5
2CSR/JYHeuMNUQQL8oeFFVVYTSOBeIrDLX8tD7bx6aAe46hGvsDB/zxZWQVAquIB
+nlcDvykHf3ub8SX0pO0CVQ6FFBjIaBMuz7xV2F+yXET6/TZU3d3wGdTGJaQNMmG
jBZYMsQ4yZ9wwcKpAuIzTecdjPMkooH4IekqG0FV5eDcI7cdMwOsfyGXWGLFOnf/
MVlG8ZvV+rxBiFYp9jELn0YmuQ6CmOyUL7UBQrvK1FN7eHU8TnYefD+roYd5t1zJ
tZr9KR0MfPh3pW2jjO9ZJSIpkl/PatQwrjJ+BdinrxIuBdZxkFjBHdrKMIcQFtw4
qFTaI/eGrlpZAYKLHwxxXzQqdSemGjhoZgLS9EaHNnR/xRBXeU7FqOHF0Iwex3eU
n5q7WfVkZ7Nn9rP/pyaNe0FBsXyu5g4xLR2d9NYAvM9xQi0VRK4R5XI8TzZ843LX
Z0qK3m/j7ng9A8VEpCO+wB8KQn4F+ZdMuVOYLV6l67QpSYsbriGl/hm9OMoXwu4Z
cflao5wOq4c+UgSfOiTxFvumAK7945bRC2wet81cdE8ASDn/OD7LJ0YY6h8/Vevz
wCKm6QlfMhQqf4OBqJ/5Q9lPbzoxHQDH+NHWfpzcr4nvGoZQnt98LUiFUE/2QXH3
ISCtS2S6vCbN0dpjMzg+k8V4XSrodx9uXqQqpIwupPFBhLnR8W7CD3AduhfcZ9Uo
JDIr8P6wa2AuLeXrGWyUxsD/6ga4zutVbPbFHnaBfl3wCp95J4hkWFD1T8Aadowq
AkkqtndgCcAhxjfgNImO8eQXnIw33xR7oj/49HKIOIRt7tPYHck19YI26EYMHxmJ
68TQ6584XSvSKrbmXsIzMdjlEK3CMHqHVhHy6wUxcW29YKKFrmlqihUbAxmwb8LJ
Tpz+dc6HDwo1d8Zc7a76cmYWil4Van6auQKf54zzlASem2qpta2VBIhraz6RyGQ6
vkFoTg8Kem44YGWRQv4o36fZBuUW1rchtc1JSvOSsIjFL9Pk7SjOCL5jovwDzAHv
nRtpICv94kbH0P/cDldLa9tD44STaVzCo3/30k6oMhhHpOIT7BUvS2+UWqXiS0CO
BxDmnpelG5A36xe2AcDRriqKqks/ZihqbwfADM3Cc4guLG3nSlVqPtTQt2fYAcXE
T1Pszjl9Dt/ThVhrFOgXxYy0Xujc3etAzngZP2TCLHcCPjSgT16qA1UxcXZ3RJrx
mg+6bJtSmvN9/FFoFoPjbUV2TobEPGAmk2FLbs0Z4rENeN2kzXGGVsLvgLhIfn8R
HA4OMzs6gghL7LjRiWutse2XTLVO7h0E6NK7k+y/tcX5hHPzJ31S4n673vl7cYXf
tyyPHBZTgtlSvJ2CLNEISirVk9K+RFVgbU7cZPeartn8g3lPs3v6XeT2n8xTSpCV
jefJ0Y06VP7sAeT/UdV4dEAtHUlnoL18WwD5M+Vwid2580kvYVdAUzV7EDSePwEv
nLb1tkJgAu5uy92+NTJDm8kWs5OgEXTvmQvXsgcdqdlCp9suZc5O29fnAMqaqIcb
hNS5HhQMD4tT5n0HONkC3QCizqOyATfgdzVCP8sgOeopypEw4GiixZpMwviSzpuD
f8FiPLDvuwdsQfD9NIyP6et92I9ebv0ftzK+LJ0WtpDbUcQqP57O09g5xoqx7ERd
7vwajpcidCsG0/sfbS/Vqww9m0EFjD7nfbBAWRyqQ+ccIlrz/WXw5v4vnMDX5iB/
wFQd1q7bVPGfnUrPG7jZmiK2XWwUK76bNoF/nx1GlZgx8XSvWm/cULgRjsLXwvwe
8W/KlS/yXIuF5SX0Rwy52NU0Dx6UcP4Hqu9Hw5Qe7UzNvnQN2NS0eOrDhdYHx2dM
9wF8VZvIBtluFV8i80nvyHUjyWLXdF0fmr9jHgcZsM0mrbsSJj5L/OsowNp0Gg2j
nVD8l9yTsW3IQFIAE3YCJ4/CKU/wi4ujdrGXZc0/k1RqqZW/xwTEtLFjXHdYFZQA
6q7kI63C0+o/TkC9l4mLFaWyi4s6loij7WcMJDMsDqSFSmOn+dchgyf3YHAvZPT/
mMTvAR/avQ9Z5QifI31c91tg+m1rNm+hofrE6jR+7E746NVO0qfEEquFTYcIJ9F3
YRmdFGUYnSWnHqG8sHJJZXjsHJ0SIkz1VwBYJxBxxXlbbL1UPoLAfxntn4gjzUQG
AFA5jm+pqDt8W6i0qzI+fu0XSOWPJiudDTxJly/cTBAX6mu+p22csaOIgqc/7fqI
jrzdKKtTG4bymH/yaRUoiwc5nVGGMHCNqyi/Rk8FpnGCd1B7QJzEDq22y9mYHuL8
Q/bsoNqQYB5VHxvGSjFN7+xUDvk8DOFahol0jK8mngXyNRgHbCz5YJnSkPTjgTKm
FOwoQgxPmvAGhwXdFQ2hmmOJm6Httjr3EizgF/hotXmQ6cNfrEUyRo5Ki3aXdjf4
s29eRshdv4eROWy5IMdhKLXlyu6GotzXa4vqAqrZUVCCp6hZ/MtZoZZeARMpz4yt
KV0M+UVXdbeho/tqNKxh4NBcsg6khSa+6rmwubjaVbfb7be7Nk1qUqC2Wu1DtAHB
afjv8I/17PQESasy3/Nf9xPCPOT+LVbecXsghC2Rwj9RmI1WrOsdntOzAmQwSi/b
zq8LnpcZFkUlPoyTJjleYjM35iDRSZrxdImUPO9RO6Hs2mvkCB5Z4vQt6TCvxACW
8X+ab7+bXHp+rFGtQZJ74GfWf/0C77WKUYsFSnDDTIcbtBuFST0T3zg090gNJAnR
OdRCjSno0gGS8KGtBxbfrmt0ibcvgJwEyKKS6mQfVgTNmLYpOrD0tmVAKb5ONfh2
NOkB6X9V1Mixr4MIPvadVHR0ncbix718lri2euSK6K0Ztdo5iZ/yUKdTF+r9i5Gk
xNGlhKJT6KAGg/Z/Z0weWtSglIyeQajXtif/ngyQb2HHujVQxjjYXYaGvficG8Yk
ZplXDJvh7sdhvXnpZP4AO+71RIpYHxO/ZUdGf/8TaIJSa7K1antS1k56Vhy7bSSy
qDV7vonwob/64QrdrOvAX3qkMrWDE+/PPL/NQ9OxmjTKlH3i0q9W+MWPeTUiqKU9
M/lX8ZRVknHyUoilUfumRUnGyZGwPpUAyxm64Ejg6/2ON4WBvYKk3zup4BCa3i62
udkqNk+cPJWIPhUZcjphLml8qUfTFAHGvqDhxCfLlB8KjMcT2HMWBPwYDoyGTBA3
+rnudHnImxsTCAThevrVx6zSmzbKF9K9KHuF34ttAr4bwrvppwZiaBRKTB6PqYTu
LbhkDw/s4oavWabWm9LdFADtUZGGmbaOt3vvJogUOcK7laF9nQ2WNb1yGkKCp9AC
lSCjglBOOCGbC9VVU8cFhlqPVIi4Qb6Bln7wCszZH8EVTVz5Tszs/dk6rq5e6biV
BsYpxpWT0GCLvsYxqD2AMPLfQJOwwOtvi0Rt34SJYKU4aZspJzmmstQ/KRMBuoAN
dSQFfoSY2tnZki/vEMj2dcZbw4iJqKNKI4iOwhWHoDRIAS+5mBxi/6rENwy4sGBr
ZhQ8DIk0MUScEpPZ5iIq6mvrt4Ipyv0i4VONfcq9rYSL03Rh57N8TJ3377kYxI37
kxefPWwh9wGSgNdgIBa3O4NU2wiJVJXAhU7sOqx3GCkN/8R4oYbyMLbvYLQoQUbu
rhXMl+mglqK9mBdnVod0IbTi5QVgHNesY/zDLbMpkQONRGHHzr2ktteBY9F6VtYt
Ud1ApwE7oR248QetVwr4MJN1tgsnX3+qhPP0iZASEOimvy0J/mYuB1tA7PWOVN3x
Boh3+oEI5VLsPwD6AZ0ElfzCsg+4nqRThOmfw+IMSs9LBiadjZGs3fdSZA3hPdOr
JofUDJKXZevObv4a8hcfJBWID1gE1m7eDPq0Bqr8XkrtEFsXHsQW6NFq/MsnwQun
sXeOpBMjNsUx65tYHR4To79zkFwyLNZ71k2vOv5YfcL2qsSBVGqNWynpFlnVCej5
vVtJADVJuOSuLXHtPNK1wH6lOoQ6NIO0kB1uD/NVnLIpC+HHlJs9UN+X5rBssH9L
qqOHpZ5GfpYqMcI66rWrQ6+rI2SnEahCQyjkYAp8T+MfFfIcNHONR97yQFTXkiAw
1b/ncT7NZ2GyyfpezoK2dvhKSOvDeoKnoNEGw7z1IEMtUbW/X4lInerz9QgjWxyS
mwZbjY26yy2HdI56abzXUg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
b6JLl80Ceis8fMp4bsc46lwXB6DG0zNimObB0GI+UVDkOVME0IRI6fF1BhJ+LJ4/
uGuki0iAvij5HJ1MFEC7CLoUidDZOsMNDNZmyJszF0m+eVI9kko3n/qroB37n6UX
G/hx52bpOlzV83VgBSfZmTdLzotdsOFbxk6YgeQBKDXxKF44HoMdnIYuHVMc8E4X
eybPOQPAfZh7SU/KNpB2eX8gzvHTZGDCMCWE0hmi+NZJABwpTnfzkBoVEgiZ9a8g
Wyx4auDtREgOBdewOQGUAHItIMlm5ac3aIFcyue6Knq8FDOtQhwwwzPbbBh0CIpo
vJpFGUkLkPtI9s3Mp5OWEQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4672 )
`pragma protect data_block
YeJvqfSgdPAccLWPhtuNWy16/ob7CQwwYLSLLwTXtc/Y4Cdzsu9dEYzA0AAajXLP
bpJRbHSPlwFwcdm31RKF/ZgpiX7dweGS64MZcRJvuiJE/j3WW+JWMjDh53ubETr0
yN6XgAgJskJIxyhVFI+rI63TTVrNdt5ekndH7k09wuu82R0kLj5GKu6lpG2lrSQQ
m4mmu6M0yG9m7YFnpgzeDe1ZY9R8w03Rw5b8234os0aYL5qlu8T6jeEHjdPdA77r
h95rKmvExk1TNOX97OxkLkr4j95qLosHkUQtomcRnOX/3TMz5D4AzTilRhyCsyqi
Y0iY48SVZUpcOUxv55p+Jikp+uF0hWNo2nVWlj/3B4xHiUGHeBgE1sWj3n5zaa7W
ASrl9YV3zs7xPA99t34KQlyCBphaAEkamWHaKiiw/Qe9JicEr8YzWeMJIuTQ7hSM
fRQ/bucFgNcuCzQo3ukIqLmHLi8Q5ZR+MdT9+F9/e+6Kxg0ulQ+Wk5PEhqYtH5ON
u+zcNO3TwloyKixjVToqs/G4kzV9wVuDVBU7odyVYLIo9u69UmuFXS8OvL3BUZP/
Yh+v8qi6HndhZ/FtV5eEwPv7NYxHo4xLA2Lo26MoX+eNDdWJPVAnfHdyjA8GdXIP
PI2XI8lf/oPIZcuaWhNuL1ukTTEn6umObwLYXQvNklXrgNPPcS7/W5Ge0sEoIdXL
DVlea21+aoSksExDhI3Lo/gtgW7GSnv16ZjXOyraiE2zz35LGBCmNTYUud+R9DtE
aU0zHMGTtohcLAD6C3iGrYfI5loQmP814i/xo8gLC5Y9F6imuQQby6/sbjaisSmE
N2QmKACdv6Vg+hLAtyd5v04xQgVC48rXEvlQe/h6L4Gjs/ssfOzgxxHUSN0NT3oc
/zfeqT9Q06oAOvkGksRQioEUgzCOabstRAs0Im/rRRMNIuI66xkmcJ5zztiUAnlz
E0FxUTX6rDKW7sHyM7PjXcT3ZMllloFOoM7bZfu+30K+cgDkNtzBGSd5z0ks7egp
OyVR3M+HZsQo+ncCcPwYzlnIZuQ514rYpMMW6bsikevFuX7PXcwgmjvNu2Kocr5r
3W2DbE5QX+bPVhrab8lHQnYW7tgdGeafJkcaJz6t6waAQv447J6YoYI0dBfk/DRI
ntqIUmn9ojOS0pTGOK0y3HWr4IQ9SVvP8abUjlT/tM5lv8wry1mIGXVZ24Sok3er
/7umO0njRIzHkrtZEI3kJTG7E1Q7qFOrT6qK59rl0NduUlizh2Iz4geisz5Dzt78
/42WP+OvpUYyWOhPzayWcp13+SfLugdYldhAnrg/OXmFKYkxOy00+C1KdBTQJTOp
5F0R03eUaamPRbNjENSnv4hYvPRyS1vlXi1m46c/FSFxEEWOBBpKMJH7F0coX3KD
2FuPLIHplTB1uKglyRsWzMZOMz/VbeNU8KtVpqWCas4KTEVeFPusioDQuiKtmSWF
dBcOU1gRdCqRiWGO1arXGGXiWflMF+gJsWM+S1l+56qbl53BxMwWDuHaMDqfiO3m
4U8sakmrIaRo3QjvyFaTEzx4dd5ikY2+P6mW4Ip/GXElBImrWU4asAflSUpzSm1a
CfZALe/X0GYeIiTSYSIzk5OImT+NDUyI+SMP/iZwHm+XI62PTCRjUKFgzZpN3UO5
Wq+EKREclQtuSsg2RZs9G9TSsVNhwf6k1272FZUOQzlrQgNPpNnqKHqSKMJgmvKb
kUb26O6ZD5yJNu6xRsaoJapT4LuMKkBzTVngeBMWOoFupZCHafpk96CMePZ9g7go
vMTa4lSvVK1Qc5Jl/yipfhCoxHRusy7oXoyVdgx3WhvkWKzOw+L2lQy3gI1VspOf
7Nzs+3lo+C4xecvsHv7SF16cVdKcuddrH/oGZPDtzBxsIS1Pfuzpb3ErNE8+EocO
Z9QVyz9nkYNe9VS+4idz+C3aTJbgyqHx+a5mNOcEkzFdlP03EQNBavDSe7ioOCH+
9nMfsl4KOXnj6ZPZIufpjV5h8vtPhZS4lI9297t8dsSm6ZxNietmuuRwL1A0YBWz
ebOYQjzaYJbUS1Kq8Y3zEx5aMpZbrd8ozxdOOFKedPLiuTvzW1PWHgzDV/WNf2sN
4BOv64LvbrUhmbNIylNVY2NosA2WVJyE1tWbywOG9J0nls3JFYCsle0O+cA2E/Z/
Z+PUskI6h2xXxGb6CpGiJnPheCWzY2FFcK4iDyTWl3Z7sZv6GmyNfhnBSqFXkt+q
CbdaANrsVPnUgEBC1WrzO/Ff7oX6yaJHYqAkCxBS+1rD+iYVncu1PvycYYgN0MPh
MW57V8hjgskVBV4XafTtIKprXhRSAhonIiKb8stVhHrMOZ87nyJKu3K/jxGFHgoV
p9Juz5EoBa/sP/CTvgWiSLyl2Z2lDvNRUUrWCCuLAHAdhnICbcRDr88cO7kaecWv
mYx0ihAwfTV3ofRuPDqejQ2jSg9l+zwOMx7LMRXEV/SvptiUu4sIVpSTrc5Enuv8
nDN9ZzNCPFrQI6xTXXgxOmdG6L9oSHP7RhxMWVxStLKEooyZpO5v5EKUUpVxEEwX
O+g31CZDfQf+MG6wiaQlw+v02yGe+1yN/JI7RKRu90RebW2GFpONLk/77DgXKfaq
dgj1DRHbhlzXZHBsZqmR0dB5uPKmMKoc156bJKppDp8g9Y35o5Q2+DfluFM6NsBl
T+t5xJ+JWBTcLj/kvC98V1VEEqYg4OPA315u/Oa8zpi9b4CeFbDeMqTjFmzre5Ut
Mx0DOI8cDBkaMGFzkwAPiHmnCs6zSTSNaXllfT4sUObGpEs6PvM/1gLtt2PiIAO2
/E2w5TFYfnEdYP9lNx1ryIsp1+WEXfMpEco7uDsCdys4lWnTawug4JFhpFAUnDD2
vWCe+3REJh3IVC3bloME+xpiI0nPiY9nRj4n8czfnSYhGhVTGnBKoPwM625jVaWM
0LXfI1P49/blm1ysMODmFoZpmHv83webXn/ttQZC2q372zq0KJms0wQVAdH8ce7D
aRGF5HD0e7QciXRmV/r8ts50lzDCWYN6WKTr/PQJQpW7gdkwWyJEyR22s6Z2Etf8
sF8DsUOKL1sf8RAruRRA9E1FRRf7W7SaJAfbfbwcqDYhr0cvPnLxR0PEyzEn/lRs
3WHDPC+p4pp//ZH2bS8ozaymODjZ3/TNI9PS47p7weean/KFqiLBA3myaF2Fd/3t
boaqtzWVEvEcMK9wcPYoCA5en6OUDHsqImPNjX69gd7Bw7FhJMPc7TYPQj7ev80l
MEs6SRfY22Nl8rpzj4tQlET2WxkXnzsfxV/0RBgd7Tdx470iOPl6WGH1yxdVBuqm
/VJt5jXpUO9ZAJxqOBLqf6zglNmTbCmwswwqzk9QV1M3mvVdkFPTOaHqUI8x+P2j
YYRDKWTB5B27sLjFTht0WOWiLoDDU2NO8yp8MGOUBXD5cqKcLrtxaPEFPcNfRCHG
2G9lMuB6l+izzIcWwQGvbz7PP6Lk8HMl7aCHz/wsCdT/Tvn8JFjqO1sd2pnsevyJ
BRCJpPqjqBwE78P/WXUgExSEgka6f2NMnkfOnhxpvDgogLU0RzAQz+OPG1j/H60t
M46HqxtmwCPHofSMFnTPWVKZ0hM+mxmBZMHu1zfAIXxQl+xKREgF2YgHEkINzINi
O7Spqc6tHLAD4JXO2FzDK3XZvh1z00iZMUZhA+HUTPxmxG8wf2eiSnhToWSI2zMC
N4vwM5qzGCF4iFvjeL+ME3cFg5X26xFbWDhG9AusfOyozWgbiXKpWo76YVSTieJi
ezRhEWkYCldIUqhGk6spChRmia/k5CDN5mlyF8BBGKrT/q2Qv5lkwPVP1AJOFAgz
95DUaVVWmTjFkQZCOycVsRw8fpBMNpbHSu/dLKFc9m2j/j924+LcWcgBYrBo4PkW
/Towfx0LGGrNld2baVZvNp3ysd8y8FQs2DzyCW1exhLwXHdEYLIQad0/RcY9ClfK
/XgruBjANW94KHdA+l6OuLI9GuCxh4Sor4H9FZ9GqZYNy+UYkcpVn8i3vzjvDJRD
w4J5HWkIbnYskzMQcoSX3c1s2mjUAVBUxP0Ukv+pVLdl0lvJhYInJW68+wrFWmZd
be0uFyMFcChSwA2UovsnXJw67UzMTOGxPe7h5A/+YPk8x1OsLCsSZy/iX4XEeR+S
ncGPl2Dw0Q4bpfQozjyoJIkGK06sJmqlajHPGT6VIjpP34k6aAYq4Nbl1dmmvswz
kCkfFgoEDNSRGB4Rnakt/a3g9JPp56EqP4oJxM8AbDJ8IEIEolKpbGKB1M/AeTeJ
D63Uq8PPCTsws4LuMS7bveyamOvSSZ7GGPnGCP7dd97rKZcx7fY8RR8wOtGjsW25
OWish8t4Blh2AikHxzSd3T1bbDRXn4yNJ255UUFtXuKbGnfzhWZm9QAZCYUep8dW
kvrywHp65drhu9nkrJWygSFIrXJOq2fqrFFrC3oB9MSCx/UF/eyZZ3VVqI/i5XdF
6SLl2N1LT/bDAJhSf9GIL4MoIMUHew7Ej9mlOp+Ox6FmGmeef03Q+aZjFg/yxYKb
CmbsmxJoPHD9ULeiy609JBrrDkBmg73bsgk1gTqiOQadJPyMnii4O4LWd6bfLaG4
wvztOomgHKoRhLBoPlv0lMKUz5nRx9//1Euc5+V//Z5ty1WZHNxUQCa3W4fbY3dv
M1rfTM8gd2R32GrOQHaZfbBWiyfuPLu8amYECaafcx6OkC2ZeCU8NKsopHa2SLI1
6W4j7/q3WvyQd0nYavlkyjhP+uDTesEbFC4OjP6CssBMwBRGgehYlmGchPUJrYc3
7EB+UjGfjgeDQ0AELBDomt6dghjUIBEBD4N84a057nWY/qV2h3+8Ep+8xhc7ULbo
PpkglxbKfanwJiie5NO8RfquK9gHFE1O3iyycU0PFE6xud/00q3KpZloRWBlfGT3
R+Ev38zMexndu+1fzutga1Kpzcpk0f7z+wqEbS/yF/1xXonlnt36WXsOyVBLIMAh
Up2EZtcCrWhnQhZaitqvK9qdK+1ju/klRn4+jPmuwK8bQRVI63DldgvVfPfLBl35
LDO98jbx0jXm61+WonRQsOl6E+4P3dBdXDF/2A7sz/t9fYtPmows8xIypBBKs9AO
QmqBQdMDSWU9XU3eo96QKiBbNK+D66iRLg5zs9kuS8G10IvOQ2kE6ICSR+ADZbAG
0dvoVL4OHw7WIHx14oX7MvKXlgesPQf6U0ynqPKdmRjxjvZIzx5zh0uvJ5m6j8sh
bMgO/gfXPnxA6YHz8pHv6CfyDu1CkdMzCi9WE9qHLTG4vzPY8p19szaXuK7JBS5j
hd6W8ph+yqUygWR0WRfr65Zive7pt+lGT7vWW/qDGUADduJsM8atZCxmqxgiz2oF
U9zibAZx8J0pFSoXtbZx6RYAUgBT9ABeiG55ym+isNZmCb0T2ViyUl4EIxjUXczD
LJTe0TVxnq9jN975HJqnFxaRJezeCjjpEhsEim82Es4uaqON73HtWIZHkCwwPnNz
rcCfGeCWObdyiTLTWYww66Mz3zZ5LM8k6Xh+iV8i0aTNqOMrUUGmv1FNMYkmlj8c
QsoBCC8UZ5nfma7iqL2upFjUXhUkKBynkzWgGAZddS6C8aEdKnwRknYxTKL15ize
Mjqwlkl2OCGwsdioN4q0M8r+mUyR9rCHG61vuQR+5oQ9+Rr4qGJiLptiVUQ+inHO
FAcn+pDJ9LKQQk92kHn3W35xWMZ2gT/EGtTNMJBqLWiOUGdnCqUueI36GoJyw4Qd
ZUBGSuh0NyTfTPCA2WG3BHQ0HYBvXloYIv8Ip+HoXGcavQXz4c+nkQ65WO+549lT
F2tIaWcd1WhCKaZKgbmolqh3fnWIOLiAHZzsU2yLQF+IlerxU/wkLYJanIbY+gaV
X+xHfh9m7f//LdxME8xCGj7zh2rtGTbHFQXxeq0iF1VdCLeLvklGO/abf6loIQFx
R93LZ18Rt0xce8alk5QXn28ZqLEnry7N8xfQFP92LGmz09YAqPeS1K7utKkOYtx1
yND2DB+8f1BGsep/l43F6Q6FmWpm+iuI+DublkXQVsn92vAL/xAcIr6JLBAOZtg/
VRpJxsfNuldjajDU5OiaN6kxVNcrx4PHg2iV7ed6DGDP1ydfqki7MoD7iRmDenXC
jeVcJZZ2GhBNJIOVzQj+K2+XWye1POZBu4PT31zURRCFBcIIfSwatNIA4wrNtgiL
MV3jbB0TYTsw0hLYYxXgkw==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
RarMbDKQ88QRycXH+xGI4Xh0wbKzDgk3O27zhW/vw3iPnJBo3AZy7JW4Qmb8vcih
J8qbW7FNlxfJtZkqR+g7sBSkURiR2k9anZdzgP0uQHWVtngXLgj72Itw/hCJS21G
zcKf3DdGi3BeYZTPoA6tIzIHCgkxlvP11QmgtsjRBKaViEWaRpmfDVLhGCdWjlFE
pFCEoFXJKWXhScGeL0NdZNogL7SGlc+XNlcPt9u1UldHbuQxMi6TeihNsEY6MlqV
JC58lUov2dP1FTV48cRggafz0wvnxtcR9BkecMFaXXeWPbKg8Z4tpelWGU7lc646
Rw4EnQRNMDAa/H2ZByDW1g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 11552 )
`pragma protect data_block
vggf9RalsTxQMgnjR6HSxlKAcf4H8RJSrFhOw9stXJW4LxKgetMp6NRN6Ho0yIcH
TDqnossRhZ2wfW+pMlwoXt5c9TWhHoe87K6cyjf636IlYJQHaNVkFNCddEywl9xl
T9vU9NAY6s5pi9frmAKxiVDhGLgrozsKtpvaqgFyr5l+vQKpX/D9ADJ3j4SuwO+9
UpIrZ6fcfju1qFA+8tjdtQJtmKCe7VOFk6Aq0/qJuJb11IFp+d9IbU7vwCKSgkLd
XvGCANs+MM553Iu/F5r5O0wPpkZ19iko4iwE9Ez4epXBB9uhTdwQijnX/MoEDfdO
nMOASvmnqyNlsZP3sEmMAMFrOXKLiG57c1rK9ZWmxsxMJrtwPVYHS9Wcvqj7kZN4
KG6w3bTLt/vEcRpYZ8re/IaeVtArFxfKfOgHrEVNA9U8GzMmxG0KNOu4zih7GU6N
ny42icu3gqJKQ5XO1LykglS2hi/WIMj6dGvQnB8PGsHfGgk3kPhB7Lxgcq10deAA
CGXE7cVuuiM6ToINf3SEzIi238ZquFLijJOaz2tjUE+MdTklMjfbxvisAJcWBQUn
oeUn0EPbi5Y9Gfint6yCtR+dg3nVHkqKEbJARL82wT2UHKsNV5GpYnOeMHPbbKU5
Hq2Qsj0TXf9eSw65pLgbKHtbJD5KyXtiw2OtfQcuZQyvsGUcgK6hFKwOo7WMHTYV
ThfNxwuNz5OFACrvzOB4AyTltizDdCfx2uRFoBtHajB1hGXQzLIbPuNouPLn6rRz
cnb9wR6u1julf0Y/HjMQA3mNKJM5aIPACO8RFDrfxSwM2qDdKbIpBuq2cMe/Snav
qwYvQbY45jCIDhaGZT30y+HLdhcwrFUiNJRe3jvJrfvPBRhwDbXyYpF2j8ZAZ00F
62L0tdkjSXK+K+1qK/Mc5Gy/QPPTwK/JIO4smX9Nr1p4xrrauEZ9gHZ34z/v1Wmz
HatHT/ZROSVdJb3VNDhrnm0LEfu0r1VzcBYvcvoSsFvODqSHTYWz/+ZLlj0gPOoX
cEgWvFJVIbG7CILr5uR/V8s7HmJYvIHSfPN96oIs/HLe7Mtg9Q3H7FN8dhUcaNJs
wYFlUEEhzAO4XUthYMuxcQaZWbBiqfGjdOrYIUz2ABiNTXAXlPmA1VFKPDRA6C3+
ebUno4UanNpA6coH9IQDwioNKQuCe9Y98G1oHxaa96lU51Vol0Kiq9JG9ld0OGzM
j3nKBbfc0SZmOekFpLJgYNNLLUv1Ot5zCyIdFI6oXRj+UQARFr7n2DwZ3eQkA0X/
apooCxuKJCNle6F4isajAANU1h1LOXruT3PmspJilhrTJDqc5dVwPT3nOR0eBplc
U1/Q5yaP+gZXwDYfXMW2PhPkGI1oDRGUm3madF4Eul0bStWhmLg4zPQnPS4uG5cg
piKlrhE9Z0ndur81vHzj1y/5RzaTib6zB8KHfP9AwE8A1QN4mQlvIdScofXTzLI3
2lHjzsqXvsBsAGiBbyW1DLMpratXjS+gGqyF83dQDGG+KS/w2kl5pGGkrCsbB+Nz
YBTMM6fBYJ/DlB63jSvWMrEeurj2bENZYWC/Z4rVG0k5Tqg245MZhx67UH3afkqo
entBM2Oyw2tjpJhDNsFSblNBEFCIvebdhQnao4hzqwa4GExqcOTtnoFyilRVAg5w
wvD5h/opzoWDrX9Oxc4V1ZFuq7CUUXUOSdeegzQ8c9tPlHpNTRSpLgUUJosJC2yu
IAaVFAVumBcYx/nIg5Lbj0EjHXL01N/Sm8Rs5KKUkxd5kwjrRSg+8bKF59jWP6Dd
jqNR78y831ocA5w0diNSpqqTtHwaldpAlXRHuI6uKGVoaFPrD0GEOGDoqm67bykM
7uaT1uIsIeUbAnYv88PO7Ns465lMulBdJ3rFXz1Y1or+WFklXe3i8qicmuxweG8f
AmrJLN7vyN+4c+TUJZCfHaN3/O70b0Q/1rgVhotz7XEJspaWm9fLMbND1fqNqsvd
o5PYfTR0KQXRe3Aj/StTtBtvtUqiMTt2uHW6KXI+xyQMFPbS1N/35SAlVb1VQQ0U
rgWDRs1OvXLgl+cfY0V1VsweVRvLDODwOg26qfPI4QqwO4lIAuVP0Z8Pk8uFyeaw
0MJs1g2J3mWEO5kvEYmBV/SePLh/TANoTdteUbLt+hNeraVSIRbjJTsHKiQmhGTO
3aMo0w7msL1sK2/9X5Jy4t0e8VFZTBEOis//oeAsjJiepRkYqMoODOsN8xH8OL9I
7cZfc3kyRzbB8PYPbcIeNykBjOlfA6/jO0vZyevgutjlnSzX1X9R0VkyFLVzT7Zu
aqD6EcZxBgwthic66h4Pm4ZK8hFxgdw8ufGKcHM2Jsn9Ua7U7fI8PS8TDVYT+KpX
YLtqClhWBH6E0D1/JZoQ0ZMUbyo/kgSVFBh/bvP3vWYRaAsaQhJzmvhtVBlZ17+j
bRfRMSpi/ifUlfuIAtn9Oa+LzZCqVBPd1oE5/vDtjmgXCSScstXc/NU5icRxJ2nJ
9ZGdJDQRARXKpbiojuUwMM/EUPSW5XOkGbZNNtHV/fqkcbWfLKOGLH+/U51HckeG
wchQ4Ofu/vccBK1Y9f4tOLZt/CzQGTGv9nFwCxOelkwg9fyIe5461VN9M24vYPKo
b2qWEs2iq8UYZ9+PRBlDWi4dIIMH13hqhuAcGrxQyImiTt4gteZvhisupFE3C+re
PYQV0GpZKkE+/wvgdrGt/G6gW7KBDH1h3MKosRAc4m6fKvWv5mgliBsBOSEFY4Yo
ffmzV1YhsgucgO1IcKv8PyYPd1SBRcETQDjoKXWG/1Wn46tx+cis7VWB3KcbxEMj
tMq66/S7bAlt3n5qLN5LiK5eBp294EyA0bwHmOY92Am2PwY/ZcqUHdVYQgwd01jX
BhXJF1UAPQHtHPhtnfFgwTx/OExR/QPAWAUem2qzeQfWXFynOVRn07Dbt3IVgIkO
UnAAr85HSi+Yw+wrVLWkJfzeoqcOzg470mvxsVT4r/9G5jN1tp3QxpLPBigHJnek
47XSHU4WvAtvWDz78nE1S3Qt4yCBfC1XgBHbobbSID5KTKHj0o96p9sVCQRpRkSk
ygflNROESmeI8RjVKiEOSH+rp7+GyoDfDShn23m1s4O4xvf/FFaosVCHMcO54/Ei
cnm6FzBRMIDMpXpNsi8j+XErTYYi2+Qtr5DN3fUlAG2QRkoGSmnHPvagx2TMNmjq
aFqI6pAUiDaMOAxf0s2CQ8RDifzzs6PhHRWPAfxu6zeg04pj1JMIKDvzOJqKKakv
8+UkcqHp1wxl3nqkw0+7hIRIvld4acJpFX83Oj1+M93cvu5hUqqwfVQvjS/5GdwJ
D00OKnJdUwINhFdox1qg6deMVFYbZ+uBxOA6kom4xtS0Lt7MiBeMX1wHw9t+7qOx
k3jKDHlDBKbnvAEgGoOiZfjKzhbTpDix6UaMMjoMv9BprOiV7LwdFv6gHVEF7cU0
ITpT9IXo7cPukzbxeYPwzA9AzYc4Ho5IRs7lv52nr6r92zVHSqVN2oBlJwBu5DEL
PPYc7rTAB1I84CCF6V+hWOKEKgOgW6gIw7FnotC5hVGml1wwlC0Kk5i59v7ijy5s
LPjgSAXC5RnNZV0BWURCrs2V+dkeknMQ7ic9KqAS7Y6JKf4ZmdhMiYuAAmpx10Xr
BSiAQUFjSFzpERP7alFrqIIlgln4qfjMloogPb3pcv9C+0jVkB+YWXdvihw5+4Yn
6iSPqpeWjDv0k74AwdtF37uDE/caeuhRsXZC5dZbo+mqeOE2WifC/zpxNXRcml3J
gkBMD4sJ/Q5K0IgdEfu/f4LBfmDEqrRFzaISgcuiDzjWk1h3ePlKLBBtJiRzREdo
1s4SNaZjCZavUMaRFxkGTDdcHL67Vuqdhx1e/5vpPcEVEaL4pZqTHWUQpI8Y4nFR
aRoFf9m0ITVROdwEYvklFT1fF6D0FdzDWMDf4L+pkxor9LJQfpnV11XkMWojj0F9
Tdo1E81YnXryWfYYjwYpUuhlGqLQ8VEdhzbPyv396uG4lDy/QeDLU3PkJ0fESzi8
/bh/4IZEHFz4tFftadwCqMNfDPiUSNI4h06pU11cgtblcKPC7hX4WIlI63KnnZfV
2B9HCvZePmEgEf0jummT+8WKFE0ooBFjDpZhTsG2kAmHBpBHVTQAVebkLkHsjWgx
cybws2bBwt878vM7y1eUezFgMCX1hpMKVRjb00H0nIzMOaWgOx6PjmdFijz1Wp4o
LWc7n7WBSYFADnPSp98BbsWKK+zZB083JZq5K0hFjHyLUx7nyGoM3NKStP5D1CvM
ovc8Bei/ya5SjC0VHVh38aaZuWCG0DamB4TiSc3UTCitPKL3TemrpOCD0y8f/JvH
RTn5Oelv87jY+GXUeKere7zZqTH6LXrLrUeR0oB43+2rVohyJ89/+KNTqkB4XmHA
sXg/84cThwFMNCX/zGGujfzpdfzz09k1PHTvG8gMVM7Byz4XMdStf/20Y1PG4Tof
oKE4osQZbQAeLWYUdgFhbfF4+I6rq+vv375zPYsNe5pAJ6dpwIo4GS+owUUaiQVK
9XvDWLCO1UxvqIRNO7LJX9IqjcJRiiGm/0orqqx/0felh9Nxp778tJXdwJMF1iAi
ITQ2q8p8Lu2x853gqk3J/g7KWno60dfhXTUn4XtJUirdl+IcuiG8EudAEHOWDLR2
k0ecUOekCnnXjc8+LRa0QIVm1zuVGn2rt76AIm2kFnUMPAnJtaANz8pnI8r6jiiM
n8oMkHefxENiWKRjEzmlUTEj6il9VsnQUrGVaoXddidyjIaGD2IEmnjjKe96T/bn
VoGJJ3M22eE1M+oZnrr8pOZR//AgSQPJgD6z31+jtZnAOe1Pj1Xnyw78aVh1I2+B
dSSx86Qhned7vi+ZZ91Rj/yiREJW8iqK+I8w6tRLmNvHQKcYDt9mX2emWicdrBbI
MOCNDO/6NYa3hH5ClAZQ+mZV2mbZktaYbarBgzndx26DSop15qGzcvd/lXFAOrjl
lh5MVPF5nFxfe4ksKeP/jGXjpp6R/3d5elU2Gc0YYmv0A03pN0JlXyMQrmvzgMK6
ESS2iglwYcTj2bGwoW18OthJHLqK73GoK0TdobuGPR029exnQUstGKgQYnksuWEd
56AoiOpTHzvDdLPijyAxT27soFM+rAmXtRcy9hjdvmC+NUmiQxTkMLiBtUbTbw3n
ozTpQ9KaiO/xL1YrSFJ5Yop1xTUp/iB4zsdoUwSkFiI7c2PW3sQcoXx9j1oDIpDQ
KlDI3Zq/5tXsxK4zxzDeiLUpLPASAH9PdgB2e2srNYdaXUYE8G07l7Lc1R+zZC49
RbRzCuDRsARgW7ZWiERK301TEm5UVfjVSGY6Qr1keoiP+vAV2AlKegGAXTc/Tyzz
0yHBS+0Z+8IS1ORaGMUFn7aF05M+T9B4DKqgR+lmdh6BfouflmpywTWbscYBb4Y4
FF5I21dcTJrakxzhfL9guAmyTTmUY7Gycs57yKW3Crd29kRps+mexsHr932vErzi
nRGIBf8uCSeohkV0yXYBb5M4YP4bXjsE5Ip/5Kj5B0RnSqcAx7uetEi2Ds75T1hU
HB6SZDmq4mG1xSu4ORncqQdCFhn2f5lhvT5fwh+ILBKLLugsS64PF5XUbbfHw05C
DrD2PBsvUx0Fl9Hq3qG2wdx6SFA0PBrdLjo3VH/lVlabYVuiqkk1yXejvQfLhfxh
t5huPftZzm/iJfrUIGcmIoJC8mretHLTp5HIlfBWZYmjKbbC7wImOE+1dEJ1lvdJ
7qwOcSkKwvUDEhX+2xACDCfI3V1X36DglkTCp0beYXjt7dw2En/bQLd702hw3qgd
7dC9bsIFOBk1k5LufzJcuWgsn6TN/yBisHaV58RPBmn26isJaqhoTmOre9wzO+tN
Z1cvoyZiufq4FqWcfbAMinuGo+KvXn5NJ0Wp1yuOPeJAp+N+Es465Ez+DuYKt1zr
gQePHNOVYK0QkSoiRUbdHzZ9+LP+VhsFGBNpgSLC4t3egUCCcPe6InVmKK6gJw0H
Tkgkxd4dja5TBDZddzXVT8zND9U/po1G+Cn+h4ONETE++spzqkjloFQJdsZCcw5q
eBxmMpuHvcWT0wVrVx1yGXXSiiC0U4PrCzvUilRxkhk7UMc+/uEwhMhc1/XTJrZf
GNN7k+57SkETujlkrsN/geqLoBoP5NRlVdMiYC8aC5AzT9RBtYevFUmolQfyAHGz
m3OUqHcbqvxd6g1L+2jU39R6DsbiJRBYvFTZPRXIqpM9X15ygXzwJwnA7RmoN1tS
eskIYK++iM3kFcsPCMjZA+7QoIt4+pZmmvUV3SHZ+qMORVipx037VxEDCnAK+yv6
V+bQnBjWpUNz+u8Cid44HoG4XbmSr8ePfBJNmC0nQx6OjcvH/NuGd0vGNIVLDG8y
X/w/x12pxhNGf7JwUjbz7CQx2AmoWOxYTapQ/DhS2J7n8Wd2PdXX1SzoL4PT6J70
ojHJRjP1jU4IL6Gx1w7J/IY75J4DOu5O01k3xugUvvCzurR5YQlI4lYs/cNmOlWT
VktlHwOsoF/k5JvVIuKxg+ScH/twkkEvBX0kAMxe+9TI0DDi9oZtsyrpUZwnQwvx
mHWhLWW/+1JQcZScGs5ghgzkwZQtebBfP+S0O/giz2Clhd5iP9MHhUwkXMfYu55z
/J/qQu4zd6A6VEO8b8naMt7rE8T9du2AdN0+Nji5Lo2WGVrRZ78nam7hlI/s+W2t
GeTWq+FuMs8YrdYgYiUQVvEjTpN0eQy+2p/lWo9ptKEP5cU+sfFSae6N3mlBLs80
kdW16kpuGWsI4WdDzz0ul1WV91UU2uANALVsQwgu5KKHXMcxce2Ad60oaMM7iR78
Euj289GhBV/EQzsBIEkNGUmtUEHfHAgZLk1UJetjLWnPhxfWLPdAWvLvwpdgsQsJ
4A9j6AnCbyL/pbp3dzo3GP254MVyQzv8KTRjj3jZPSm8g0I19uVYaGJtx/lmKDeB
FERqyjKX/bGndbla16kg7ktxSh4/2Ob5v+iMK3n2/Dkwy0T4fWleGekfRhE/cdvN
FMZJT7tGUb0bHY8SYN2xWi/tpMJWzORejQsWZv/prD7aIewGmwQxGlROA0TQG/L8
TRFAR+EaOG9uDWKWk+9xjb6x/quluvQ6uFBMcUv0ART/N5o1b3DRLAZNFAlqn8MN
Zrt7sbGQQHzDjLZ8Vbk8iCkp1DQvxqzwtDFZyl9pd2h/PIUE/jALjQKdMo61/wNI
7NiViGGr9MCgv2hyhmLZkZjDxAUug31G/mgN9FaUk1GySyQRaZyACF+WueCyJNZc
93MW02pf7EicDvNU6W+kj9sulYqXKFXsiMLnPtyLE1/wfVM7E1u332TUXfg25rYS
K9yFN1CTsZ7QdJmJ41tzfrCvjrjq38cSxBj0e3EYCagzXoMqu6bGGoOwtm4r9O85
Rsg5gCQJDy174AqCMPrQftsjUe0WD1bM0DzvYXSKCCboBvI85yUsVvGoi0bJS6kA
w2W8aQbdbjc/+2QjdMoRnO2KJEp7KA7g2XSrGbl18vng0RmqTiXuK4QlHRdHrolz
bEjNCYinakZ4KhqjMznYfjWAHGcNjGbmq+8ilBWY0QQfdRPbUxXv0hL2wcTSwLdL
q4Wtbf3v740IBafG8Z9JfSJTK2B3bFaS9xGWQbvZP5lCDudRFiSiL1pwjAzkMr2N
252QCxid1QA9NCt3Fq8NhDyYFbzIl73U5hih4c0KvMDQt4MXOPqE6P/5S8yh/K7s
rb71Ir6XeilH6XWVuzkx+eHMyoEmTT0EU6OqHTkGBVFabdVq4gyVN5cVEBHYza9K
192o44QYT0g2SAqgSpl6sns124fF7dztcDdjYvfwvEWrn7WPas49gtvqrLcPNZKe
Kggxtpzw/62SZgZfhHBkSgv2F6ZZUOuwZAqU4z2hOYXF87Z+Ac81YS2Uq21nyHTA
HwwZVhWC7yxJXfTqiYd1doS67cZsjdMLwuqtR0tGgymMdQdIsLKjWDdYrbaT0BbL
v+98FPhsuWvCdQe+M6BC72kwnfhLJK72Uv6UOfxD7ycIW6Vuak1YlR4SZeP9hZsf
4TTv41A5SZFCSiYRGTCY36AAc8fmpS4Ma874RV3dmEcbxZfgKBCYVF9i/TpsXiOF
UznoZWw0+LVuFCfdMfns8nuuzYJw8/neR63zOf0busxpNQfVLnNxlR8Uq6jJu7rZ
xz1Kt3jKAF0rIo2EHyUQkno1CUaHjX0KgGK6ujegOfPdpC+JID4YvlTw9Jpcs5sH
9jc0939UAvIjIvpl6qPF18e4nSnOQmJoEP8H7lPpAHrc+DfcWdDxkzg/VjDNpEpv
ymJcjOlY1HM2oLrCT5Q++FYxE8brSDbCYcJTvJgH7BOfG4tTBRY2q4l0iNbU7/+x
jH1ttPKzEqKNKTuOFeq3Etsh6Jazvi9bjg+1qe4iZaTIJyW15iOH5uuR+LeYw4wF
ubZy5hhNVzXjIcmVCdTG1ryVYJZ5Z9kAf0ljxiLvWJzuRGmwt6YE4U9/IhHZQzKe
JivyFJRMILXm5dllTKRJMKGVgDvTeXD31a29dOcVz9qqv7zKxqQCOXGA5INWY73D
U7NdhZBPfTbAWH3tnrS8dlAxkg8117cCCo1yMxincFr4Ot532VMMXD93xK0pY+ML
n2CBcYwiCfNHky9Rv9oukYwwjgf/5sIjrn2SwYH4QsuC07Jn7neiDp8eOqN/VEbi
OLm320OVMzjvq/KK7PrhBN7Bs4db4F9LHMmpcfN+1HH5OQQs5VTaZJ7f2VKwTmah
SA7xCZPP7LkZcB9K1agzA+OUqNR8+38uVojdLAozHEAN1PAP0uCn9NJpNZXcwgOa
J9AWtSrThZVqfhL1AM78P8Y9HiM9nEJJTG/JY3mlcXQD2XnWSLLehpVuJ9XZtWx2
mvPtho6+4FKMIWNPwP0QMzDdWFPHcSDZVTmj2EelIt/E0d34czFLEc3/jfyx6HD1
gyla0W5/lh4gkP04fB9L7BhUFT/MWacuISwprr7//H19X8jLVku9/Yi5YJYy5yVe
d4DCVyqdfBEO8D/bPL40qR0xX9HUC+5qnHnc2T1b5Z7Dv8ZX1TfHytITEk4AiKj2
qPkboZjZgoAlk0jfTLwckwYH3XqSHWiLVS/9kVF+xmD5A4trjN5QakOMpfrj+ZbN
MSHWqrULObnlvIggjuewhIp77Q0tDpp/oNYRXDp+3edwOoFQMNQPq0XT774VYUDh
KtMcXpVH/l5TNAiFPptWushe1V/N9hy7HBmbDxITaOJZrg44kYs50LK0DiRgg/1R
tNVonB/UUSjZOJIvZ9c5S7yFYUCbqT/hcYkOFFEkPY0M+dpUq5UY9DdE5Ef5yiZl
ilgpV9R8FDEmH9/1Q0Xno/BwqmuSh7rXbMg2RinXMqQaFaK9SBb5Ci1f+VynlFt7
nE04/9SyPoOIXB7q2tTHGn4I89I1mgtwZTnn8vdMaBH5UHFE8ocfIJCvspsZqew/
PhB7dNxM2SRNL6AnodXddMdFMwMYSoZw/JNWjywjB8WfPh7fPifBvwh8ePly8UNA
n/Pn/sEMkbZSYwV9WlpVcDsXcMUOmlH0jwCckGquqkoXGJhBrpLn0O8p5ykMvqVP
gdjwRmF0GOMvj2THv8Cm6IWrnFLgl81UIicyHv276py4vsIoGXmilJ7hnqHVMHxF
xNCIn2qwGz3IiZo0CQuCag2E+I6NC88nl/j7ApdBKigeECTEk+C3wPINbmQbHXDk
BMfdF+5xM8P0Sp9E6xxiUmOlZB3SiimhVrPGD/nFuGMgd9HfW/uHK99vdPWUru1t
7X3YZpItfbCWk9Vm80+nZp9SH/bFtgDXfGKxtavlPRKswReTvpwNpBylwiBWGrdN
FNBMjAP+qODoUfnpKCI0irnauBDHfr4W8kmTKiXbkf73P/mec1M7A1ihUVTXXEIK
VONAWow6TuwKiwAFUvIKjL/uzJhFU21Zp/KdhOKV6cpdBOfbGzRdmlIAWqMFPuDU
RaLaareZBCMu7VcxtHJH3XIn62LVx3j64Rt6JO0v9fohEtQnJnRRS3hfhX6jfg3W
VVe4HC5/nnh/PAH4aKsJa8bv2ToxpAIO9doZ/iGjjhpz1KUDNx99B4jFC+Fc9IJC
QwVBs9ts/j/1C+WbDB4VqVxQrhgvMjB61EFxhd+/X0IhIPBQJ3dlz4tpaF0Oesea
hTZIbUWTmfJjN4sXvaoYa+A1M6vtEK6/kctXfBHwRhCWQNVmUS6BeYm+In7/Rvn+
WElKdGHb0q3NOq1olSUowE4rpfcbVjpx9ltVVGkJCXH/+NN0tvTHLe5X2AgiJXGc
KxGXup0BGCwu/Bg/YolTuDacKLJmZhM+2S1G+CQOmCgX2stC81Xg16xDyEEmWR9x
0doeGMrUKiMT3J8QxhWOfod21U3LfBk0RuesOt88CSMFnAyDIYhIEPOh/UI5B1KP
LLEznHLeE6LtfNKyFK/NiDYek2QjoA38V3XReevtg/Bdlh/MTHOTyHmPsJLwQcMG
DJXUEqgNJAeFXh5iKH0SWMgS2dHLRSOr3lV9UQpDw+7CKscSWtzMq9UXhQEf/OLZ
UE19YdmAV3/hzZGgDWArn0Yj7I5chpLPefP2jM92Y7J3d3OLDoDf7la2+9Q5546J
YeyCqSdv0K9MnBKcEsJ1roBlJp5TeNUq2oFSjI4RFEXMJkVYqwvooZgHG0W10ojd
Bhff7Oql6czNZdV0EYDC0KfHu3VpAvqqMeF3EOKv5En9ao7FnqI9wd2uKxQGLtLO
PGGjTQgGmg+UgshAXVJcPYobm965Mr9iprsTGJEiTi5yRcIKUWGd+Mf/p9bBSXI9
DdmiKXx9CzQ0w5OYMjuvvxbVwMmO1tYYsFYcFm5xyjIT5WeNa8kb1S8YWuZop+K0
CujaPIPqc42YG1EP4fsozW9cTUHYOO+zqKWGIifQCrpuirmVEdq02m7dPgNA7cPb
GLqpoUD6M+gGjNnBSdH4/VK520j3Xt8HMdsovXhy4je8/L0k6Igtipjo0D9NM9we
8BCMXJ4Uek2dLFcsCmkBJcO0fO4/BSmEmEdEvQZQ5A0n4dPSjb7H2O41X2RfTpF0
kdJxY9cqwUp20MO9h+755vYakk4y+Ix+2FTRXutSOgCfimZC72rLxLKd4zGO4qZe
9gMAPfYoGGvKmNOlnDQl5T+1DUYBWTf9qi2ZOSCYpBVOOHbxkByf8kDoK3tHcJsZ
+gu/2DfrZ48b8XnputMoH423AGi4Q5UK/vDOpnIIwO11jYy2tlxf3Humnqmd3Lrb
/MLQmQLR3231brtECxoQ2R7CEtnerSueyDiuKJ8AF/qFd1pRWXlJK4r/ifKfREZo
cdY2d7qUYxC924rSKjsr6uTG+gMfgThonRVju9GYaK765QP0piBct1OHRg/PVXFM
jnKOromVcJMzXBNGHWxSihzOCvFPu7XCbnIxEtoo2979+A6Bttdakuj53FvuvKTZ
t0Ru226yL4cqw2jnZioOgeF7e4KjFNmibzvSbV512Se1R2CwipYcamjmGPirVXr0
g4F59csHB6gj9jbL/2fRBCoCuM5/orm7KKvEbwQUMcvH016hlkyUQFNFgXYAz1RL
PculAHrXiCfAByM/P7EOF2911ewZO09LB4yt0/w6MYkwIykzuvkriIWGGWcZ1xns
9uTz3ZbIzjignHxhuPEiIl1+niP1mlVVjvSd8Ja7X7NFhBfAWPTs/mDscdgBV/5u
Ju/tjSgz56SK9Q+z/P9ljrP65Om5s50xwQgQyi6g82u3Y5fCxdAWh6/KcicWUNLt
iNFUJANfuG/N/mj2JP8g85ve6XpcCpuTgLoLGNwRkGJo6yr4QDget/iuow/kOxSw
7TcmAtTLtss3AXOSF+Zw5jkjC6RUvR5SV1zRiK7eYFFWWAhXjKFbRDPD+CBCaPyr
otskwFLiZ8wWIiqU6WdSgmiS/SSC0WvkmwD4mmxIj/td/bdC8cgg5HYicIoEvgN6
BhCOQf7kUqtlCpD/EiCOEfu2Jy3/1GyvIBVFsJTThjCy4HVSZnMZbnCt8r5HyIoa
yA+8qd7JQ+L8fDOJub4ljGm+klJuSYokP33eqVF3IL5pqTUY/kQlyE5wxQI/bZ3w
91De4D3LJmJgxSsSsGI6OFqefP+48sbxhjxumTlbWlnkUMP5EDWAWRNRZ0uSXNLr
otTD9jde4nBSEXOPfQXi3itzZq6GORTsC+rp3Ox4wxFwDBnFg7Lh8wE1+TP9eA20
w607a4dMJAuX8ILg/PP7FO3Ki4tX8EluP+GRoWmWPIJEOemKDX3uUqf0ddrxZH3L
Jr92iG1onTQin/pT/6VXrnm54MNq+W4jq5AgAiZ41/Mo2bOvDyfGwmHOZb3iriVE
35r1wD7HpF7ms8v8f8w9M0GEyLg1ji0DUzbKuareeK9GiurJSkSAXNlQc+IJzP5t
2R90Ac+wX2aUN5UsstuykAOg/ETJvyaMgq5vEY0xlQQK5w1zhTjor7vj4Tkj4QLu
B6qDPnBUJmJYTveWMvi3HRYGdUi71W0sICGSK/56FeQ4z///I5WxSEtW1pF1nCSK
bchfq6GgFDETb8WM/nJPbnNju84NH9j2XHmLjHcUWXSDXSWILL3ndcCpv1lkumVJ
Pc92z3DUIWji1IRN94/Es6P4ZSjM0ObNIlEClgtU85MosRQSahQm0Hbw8eBG+3qn
VMre+F+fVdlTLUScXZtsNIvTosSNgfSPgqputYcJnOGcMgRzDe24LXcARlNa1np+
TBVWxwjTHBD9KxePnbqZVucHfMxQ2q1hp9+lGmC8AXPQUX+dWjy8GgxDzTMZByCZ
ziKEau5XCLsODFmbJQKjVwn9JGRbik+kMvx74ut3FI4MLlrEgyP0gX/y9u8tivs5
nWicBiOyMW7LD/TYtoJ0vpUaA6nSBid0TWIJoRN5ygxULTZZmlJzaJKdHRvrnMbi
2rDN3OysPZ5OX8W/djzaYOWPnuYsx+Dmj5dU608eIVEe8MEbpc/hIIc7jr21jVLy
q657SvmroK9b5IV/Uzy9/lrJ14bu7GF/BNA8fMmqMwt/yEBhnMEk51wrwpWjApJJ
ljj7Y1J8jF7gQju5fwRoE+ScYqwSr8hlE67q3TbGYlDdDUUACVsANTGK0RrQWYiU
vWF2K6PkY8iLW1sHqx6MB+QGljG94UwmIXKMSUEgZ5ah81jkPy0yb5z8mZpVkrcC
Y2lCpSoClyuWBSTEmUR3dIGf59p+QWzZEmzNnqVPVNDvDwH1x6chGBxXXCN33VqO
0+bupMIILth60km5CAvuyC4q3MZJxQ2VOuYjpeXdMqVSaKmqufUgz48aQvyR9f9/
h4NMVKbdGCxFgLDfSdDjbkM8mzMiAdSGlnI54WoQiT1kZ8BGnd7+xrxl+Gh1lJcC
2H7qtnRKhmNlAkaFky4Nj9B3GxfuTwl09facgGkE3BHOuEvSp1NbTqVGorDmq/9y
GwjZM4Cdpnb6J7NjAWZvd7q5fpMaSPbiT9tMpcCnTJmq7/4lo8/9tnCeBlF//CFO
hO32uCnyspog0K4IQm4kuFfnHxRduwh922GaD3wN0LfuqXPh0eWKcKq1FuWnrR7Z
3qqlIVV8GjD8Doio+tRJYg70lkJOcbG/fxka9O4unRRYYnn+FKe+lDKtYpO56HKG
zTgYgDyrPsmcgOG7RpZ7MF/f0gkDc6V0cD8WR2wkgGsqqS5PaTD70yEmDco9TePs
BRYX0w7N/mV5Gxhjjrs7uOcQcCbRGZPM1DeUzXdQR8zWZRmHNItsSd2LXqkngecG
al/jhL0gJnU+TXXk8AN447wGzGsJI7LXJ+Qx9RzC43q/g1pqDcjbVQSPljuX7keb
kQgYRsNDsYzSUjTGMms7FPLe4nyxUL0vPYorNNtYcdJnDb+hZ4Oh6XYKOV+H8YWb
qMHaAFZn3FtUO4MlhBVL9dQJAups7u1rTd9qGP9gAieLdVWsPKuiqGYYc6PJFLn/
94+sSlslje0gu1QmpitGjHbSg3vwbFcFERQQ+SKpnVXOhYPK0N4YCHDZ48jgZoG6
hazZqXLar4ictVBBaaV+dIVzAjgqWAdRpf/PnhWRdDCoR3J4nyY2NSG39vS+IO8t
bsntAeXGdRIdzyKKUTEloNGdA18E1T36LlbVW1mJLAz6bVP30rpGuBJBZo7k2cOQ
n9rKPgnJoJ0FN9jRw9vDlAJaxTDpht0nDbOX2w1shnFAyOkR/KFAVeH1lHEbZOOc
E6iJm2fknA6W8N/EA6OE7GA1xm6CYhCin0gYYgOEUyKxY+ZAl3KyfqtJW5izJqEk
fWjOqHWORfG9/fPGODxoKsDip2cew441q727tyhYXPQgUrT84vsiS1/HXXUsWQfv
fI2ISoZF2Vj2kJiSrDma8bG+/JZ7JHeO81uoq++Eo8qYK/fqobBnmNWIVxXuxZkZ
K2QbPhnoKbWcYU3RtgoT/ulpg40hxP+7H4COGjWoGLFHWZWZn7nxD+JlzBg1Wfb+
z7o4C0d0tvywIwjK8BqxKRWR8qyq/D+YOL43PIUO4kupRUdmJ//BwOvlXS7PHfrG
IZAeNByFDD8k5JadWaJQkU6OeYX+AESnvrJxh2UNesAA/V49er1rYAP7ARa69N2Q
G0vdsGFZDhDxVObAgqsA0fuqVcKtltOh1jAugc8ra/xZ2MSrUGHsW4yjBcCSd88K
Pr8wwJKm+Zaaw1Cs8BBPYXa6fARTxaeswv1EXc+MiYsuuuQRVLRNPJLsn6a55rJB
A2p57TMcUcZxLt9iI2FJhGaAdnLjpcAY60nLvilokavBErDWV52TjQrD8T5+IImr
M5SNDR2yfBAaoTkD7eC3Z1oG9+Up5xj0meIHThixi+4U3YvYpJzrxlXnNGjjvBVA
ZtijniWVbm4Otmc0phlZeGEDbXkhG+bQo13B0q47aymiFeOLHDWtABfQ31nB2gMI
mKQc5jEudOixZ3BNmDio9yGO+zU05dNOBWHRbt8jX6s1jnQ2wj9t6B8tXVEPbvIH
bTHQhipBfcg49Yj9pngP6etUmhr19hOj42PWDM2fmoZIj8bOaAx+u+E363beqFRL
YqrtbeH4ITfD3YBPC5zlBmLoyynycAq2ZjjQUtNyJe1aYgCWkpdLonIlcThJ8koX
MfagIwS3bddhO06utiIl9JUXCvfCzgOen31wJazBOCJ6TzbvCpLr5A5UxznDBRnI
TjWRC+G2ymasT1n70c4hGc8qsVFS/UdLmFvau0z+uJUeJbVc76CNO53sK3g6t0dK
kghvZXDPpHVVLf45/kAUYUg6Oxt+Se/vOUytQiWPY8fn2hmJMx/HZn3XXYuh6wmM
4rTV6tikdINIi9fn2YR/eEs0GlSOLfJio/Gz05Ro/MFmMUoukPtgYefk84pOgdwZ
qtr5IA5CmxR2WkrU9fQtiFSOB0yC9/qjPhP5RthR4PU=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
D5z03yNhOojc2yxA0APT9nU80Yi9VSZHzyVhSdkmB1bJXsbTKzXn7woKZtEQutbI
s7T6Z+Br9ciukWFbvt2AZz9yfAIbPzKd83IV286yCTtEi956s60FHjTmvOOZgJ9R
Lo6eeJJuxv9b72owZNPWr+EKZuevS4MIUQ2k/eHzdpakZOX3eUlaXLReKW2sERtw
PDnKPX4oKcAJFpR7r/lVfCEIiccWPhXfH8sIBT5vfxSH84kjbxtvCsURs2T2y1C0
EKsGNdkznJFpQ3BBH+SbkiwCgTgG7E/luXMuYHmstn3OXzzccr2uZNm8p8tV2QKs
8nCpo+oRDOT0iIERrGfN3g==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 31312 )
`pragma protect data_block
/Q9nFCLu9CjJgVQSRxRXPVu342PJdnA6/Uf+qA4iwgwNTbFntgw2rZPPGRVWXWjh
2t7y1P2B18gkgPCOryzPgBl3yTjzG72vjZXXHh3Tric9LT98KQFk0Y3+oSI+lVAY
lhKeCgewl2MEs/hqwfRR0EUkH2q62Tr8DARm5ousJBbMrfebM5nAS5wS6qY57dtZ
IYis1OneEBxqTPU4xbv/37lj2XRF9n3FQkycPPqGQsuJuGn8NHyIzyvhtMd5GFj0
XmtYimVNk6UNGRtKspgT6qtFm9lS7i6wvhNzpgi9wONEuZJ7YceKj4SwT4UogSRn
Gnqc277YxnckCuzh4cdDh1kfXE2uOBDbdayGGFoRwiOzTvgS9NGG0vnde18Yt4G6
B/5C8yu2y8PP087IIekVtUjGEqdnchdYegpN4hRJ3+L3bVt2/oJaX141sjAtM6ZA
xVhUTY2IxDgnex2+L0DIbdYq3sx2pxj/HeV5ZMD0YNm9kBQCB8VB0HG+fZCgqkVO
sRYRGana+1X1B4YHX7J3vGwuDdLsDH5ac6ZI148aB9r99O0ISKQBUuftgcO7JeoP
9A/gpJHFJGNIqx38iw3CW0U2+zforEjyrppoNDnUmSggaUbsTCXIy1q4P8TiUkkZ
xYUVne3F7VjGXK5V/a0Ah1mRgkh0cjtDft9E8CzsoxBRhwmEal6lZk2kEB4lUkuZ
+lnFRa/AOZ3E2VHDkCnpcWDsX+YsVtQqdu502djykDeiuaqafZGxANh5PEypmTmK
484APTNYIxQByq/HSsCkAjaHo6eMd9H+ptJoxsfjtdH0ZvjrbQEywG+WRbhplyRI
7/efQvEb/AM9lFd3huMkq3e3B4vZYaVVOMRKgFfBN62sSJsY5WgqrfrQHwCwJesG
qR/zSMusomRWcjmO+UqIG1ktJuILnEnv49AoNhnwzwmfTUOfhSa7nrKiuxiCGEta
h6D1nzkKvCRPcCysWL+Wx58ZcULdNBi2IbYPXFSWJJmFJkbgnSCahHHoAEACxzyk
qkAhFyq7SYLPPO46uG0pSpPDImcsCTHW3NZTPW8aq2C66OlCn7VwZhp6AI3EgU79
ByWkzAJ8LlKv0wNoep6wxe827nWuEmDP+2l5ESY/wclGPBCojmhoMJ9Ii7+lakNZ
PlpvSMza/xtoI/DWzIhYhQsGfYohgd2VRO8QUdm4I5zANDw8adSyygaqO9o2BDWK
laQH3Ur/iL3+nOKc16nRKovUG5H+58HfbbgCeSASRPwuWFD6J6uvnhPXLT54SG/I
QJMlxj26+mFJzGMGwzgYMRrBIF/8lakHXm+jayEjkbNy6d9UXMFkdC0bCttRt6Z2
q/hF5VprVBotRYtDjTDMGLzY4KTs9avnI3IIbzzrYjZbL3PtFpa2a7ol1zD6r1gn
KBMLzKXxbcGUIZq0gKEgsT+e8G1hCae/jzEn1PHP1Zw/GEOtDM90czggEcCcxDH6
6UOwYt8TgzHT3hSmMifqxd5rrKlYHVj6gN2L+LW1KZnxbH1CsvKa18IC5bXmnk5t
dKwMap+/ayBLnWmJjjpuZchA5w2UXGN98ty3jnxao48RfcAf8IJQcq17N6jv+WU0
dpGRvPWnumwnYAZVHe1D7KUhDNrg16QVrJ7EB3VpGbjsL9na+RtalGbLoqxvl1ab
28g64EJuyJE7TjiYeU3MDSE7tdwAFGthm0wVnNRNo5AUbANMHHMlUW75plad516i
0jHwQZ7K55T+2NEmxirBM2p+L2OTF9XGcUSWdHn5o5MZ7xLMW2HYR2u0T2zus7zy
kaP+480nrX6naXULlDO2AvIkikDlGHojticlLEEpxyZDiR2F9jYLDud6ACRQwgyk
urEK9hqVTt9+KZYqj+CjZMN1+iDnccHagJPnTK+dNcMRzx6QLV77JWadCIXEV6Jj
zjicrqBxQBxuFwS4+LQdFPkVjIRXn1kmrCnmiANEwrwwz23bWptByFcQOtkg7sXF
mbM08ByI0ZZuntvlOEiq3U7rgk1gX+HmmqM1izWWRLwQqy4bUfNjO6wKN0yNr5xV
qeTW4IAgj6e7G6GeCPDUo1XBaLwgKgpaAl7rFRYfqWMkg2b645eB65u2qchNzuwj
QI4QmBpA3i2tYEGkmO5NaYPNtoz0R8J/15nRCQMzU+bnmfyZLojUSX5HMip7Rfgr
oR7hJGN0si3N4K+Id+i67+wFiSQXXbJetJeUfBv8g1W+ZhkK9t2OV4ksqPdUFlhQ
ZeZtohYjK3/4LHpoz7LZs3wPCBm5dztXBUns1vgBqygIR4SsJLbCI6CSLAW70wF9
UbLTHfnyO5ycRl3qcJLBVuZ8s4QEXkCNotti5sUAMsSX2qgstBKcodVUcRI8IvCm
eKLs9NmV87qQiCMi0fRhL4jx84fSXnPHb9i0VWox2ax2WQpevl0kjpMuizXvTvhP
N+550bJIjd/3mSEMiapWK7Vj5lwd+V+UMlQkgVggEaxlkrgz1DxMgkctXBtsXzYa
DKCxOCuRWOiPtJnL8NRRQr1M58e8nUBYpz6sjfxR9DK9HP9FFenu+EJOH/Vft6lT
gRkx8JWj8Gqvd6W+wC7hOgUHxODfyLQwOfxufornsXmL4RzIhnlC44mFzETZuENf
ZKs+ybs/c63kA7VHad/BWjS9ltMc1t9GqM50sG4VugFZU7fUfUY97TUue3zOpF3y
cCxJnyOjI7uMJoe4zsSNE4CR4tcsP9NMcCcSGOp/WiXklAgGWNpGDwCyghO4kSTr
812xtuuYi5ELfVUmpOshsY0UC03mciiIJqUEe9OLoT+Is8xPvLJ+3O/5TlBII3K2
wlMV5jMt7nKYY3ftXvRoxmuN4oVS7jcaT5E9nOYxzs9Mwqbyi9Ye450lVgbGMCh4
oLRs55Q94t/+pp+RV1BcbjzkumfSp9lDsQQRr+EbtY8Y9hZWj+/MAuOSLnvUmSbA
YCWnAAom6WwFMFnLZxKtTSlZGnC8PiQfNsbhcPTdzI+tfutM1J1MYFC5USd9PMUX
vaN2njuJULL7eYs3onm6ZcCnDDSFX5xAWjEh9u/BHOTnRKnBpjsi/uKG5HNL+p3R
KIr8g97bQGYBAwnHNkVa2u+n3dTlJcX58z/cfDXpvB5m1tcS5otesEBs9aYK+9wx
PposVrO8ZvL35K71Nrgi0TY+D+9V1Lp4zZUt4GXqN7zh0srqpvKBKuwZyy+YVBv3
dK8QQODGl3t3mon8CFrjAo3cNMTe7g+BJ6DNIYGOYGXg5Pi2hxAWiw+G4C1SveZ0
3lAUEuG343hTpTWY8jrwIockVSqUYo1VJAnF7gNcyKR9OT7CkVZOGJy2ZsHSzcvc
axzcFGu6o627VOvDPiaF2aLvUxqVkZFgYbSXK2wTM8KycOiyDABJ18dtjvHEc+Wd
9zfftUfEFjLMW/AWRfayQoGUgMUyRHwwrRTwomvZDaEIH3s8ebx/F51HcFOXtJhH
2/odsBGGXj8YmaosBGyFJgy2TyqEuRDBh/8Atrf18Q/BnBuzy1mhobgbYpXrqPF9
O2/czzrCSm/hQwBTpmgdcxPyHEj0XKjLqYHrAaBQeoi0YiAfzIpIZyn8IAGflM3X
uhHmAzrEh+xbPsKarnfuG14ElR4iikJj+sK5WZ0XpJlupWaGQ4yGl5G4/Ai3WR6+
QBnVYpwMMzEmG62r//UIObuLk9+Mdc0Um7U2Pom/c+iv1lmMGcZYH1QWPi2v+6/B
uf8B3X1nf6w+7dEYAGr9/FOpYyUNBg0Yc/BcO3u2pOzDWV2j0O1NdKFgsGVCEqgQ
f55Ps7UoyR7HwkXjdlcahm0/VDcT5YAaciW67F/K26vlanPVZ/B752Y3PNCWo4fA
yRJZC3ZdGTEnT0u2G/3F98AKfQV5IHsudu9Lqd2nVHSSjgb/PIhCnv8ATAOYfx7u
wiUcDGDNCcrZS3pD2o5z70iu0ZvtwgZA4Bqj0MucREiC+jz373L/NaA8lWehOYmj
syE8Yqz59VAJxJ2fuFbcGTHHXN/n8mL3Op8bg3SURhQ56x1tOxszOMyXDmlXPm5e
sPCmIpbN+emXeEkJu9WQu+q6Lr1mZc87vYliD7QMooT+E6ocqEmzTkpmgbghpYg/
2f+0Ig+TYUdyOdG0lRSAn1WmlqUCHW1Pel1Nj6kO1XoZCWkTWgezUtD/UFPMRZZa
mNO92OcF8iFmOfBlpAeRdN93inAqkgaFxGbd3ve9US1XVYmHMJJcVrpZmCWcHX++
dayYfCnVN3jjdCtu56yqA4v4qoWpVjOP72I6fx2B98FWiIRNU4eScxENILvq01SR
+/jjV52jUpMKaFAXwFoGvYUvpiWzdWRsEkq4cM0Lfe110Gzedpbqj2fJvDXiKD+U
4yu52sgMrP5Sbf7AuZgdao46pHtxQauoEOgS5YNTOyLew4eqdnQKlKeYLDMZK8hh
ZVw6mjMtGjwbRHoda0/ctaKkiqBZpG6dNw8QSjZfSdAmvzOr/TKeeuzvW3AotwPz
9Cw4sBYb5LMq/IXPBJUi9KTu1ppEaW4yweRntU6EkQlHqDiM9GFxPx99HjtJmT+8
T68Gp68SxI4a4PdnZjxavv9WNK2Jj6X2cF9spyRVZiZsRLz9XlPPXxhLJaIUWwrb
zzj74l1NAQ7d5RRNGP7oLsL4/lPB2zY36j1sPiMDNVhOCQbWwiKxcmAIzBXntDS5
ssBSJsJCd5X2r4DDGt/r0Yo/zU2ReYSg5Agi4iQ3DSIYo3L/sjInqoRFumz3xAo7
17Ubm9FF/DK8Rjc1Uldo51UU5qVADlkSl2mdvJGjgyPde8N2Vqz+K7Kk2YvoyE5X
CYen8uMN0B1637ZvqX8o8JnQyYq+9tivXSAvCDfoJSt/eFiFHep0wDnEgbjeF9pw
DjbcVZrq6hMcvLtSCHZQiZL3ZZoVSBZJmKeIFC+ZO1aNYzLv8XhNRBQkrYf3nn0w
EjFmoGVmseuEDdlXsf9mrabdPktZQxT0Qphkn1X4N9nA/jAYmL5DAEh6OKCCglgn
Vr76XDfJpT3T+2IOb8SCt8qT1ULBiTtB53p33U77+zu6ApD4RF7idQADsYxHGOGl
0IrNw1SUlxrHd+nOH+64WDfb3SRD6b0Ky89+w+7wfaHiNLzkTtVyImXMzwbtMSbx
MCuDUV8PwAllbWJeOJHQRcmooXTQx31rql35oUbFLsMlguF+3dl28LvoLmHq31Yr
ky3VtRZv66iTWPzz5rT/2HTs0GQzloO1vlFeIUMUHnRMIrkWnvYCh8nJ+4HMXPxj
nTFFNLSR5R5w9lwxNesDqJ0rGpGyTfXawU5hYcQJOGsk96NiuXSjJFGM0s26U1To
fZAehT4fOtGjiMZ01fLcE22OBHQRxyAA4w3KKY4WcXKbv/TzAcTtkj6l8/0TC3ym
irA7zJpMi4ICO3yHJXPUL75K9hvHGKE1tKrkIsR/jDvOuUSXSiFoJjulNRIaD924
onEdBJvPtj6UtIbMjM4hcO37ZkAYZqioVUjduHQylqi2Bzozogr3nNU3N8bR/jgR
4Ylwh5UYyEbBp2DqJuCnJdCo45ISj1kyMC7aviY/M33ASSpxToa5fiuXzg+ZnoAV
NjEtbHgIjTRYQmDNerQ+QDC4GOcve1IhUIE/Jv8T3IFY6WhPjpCV55fkb/SvLAe3
9dlyN5ODSH6zHYtVowhbOG5A80YCRZ5Vp+d/jOEyCgXFTPRNLSKwaDX8SkMYyO8r
d6X73kisArU2GaObot7Vgrj6SDQ9Jjv3eMGN+DGNCo2YZazayclL2Z7Uo/BZqUP9
eAAtR0OZOkdbm/edium69imQRDaKJfHRQhpO2/4CJ0tBFVtCi85PEM4dIekxSZdt
sO7Io6UeQhMx5UD7DuX97Mvvb3Ao6rIvS7PkQqlEINzNq0pGunvxK+kfPgBzEZxE
3mGuRL94sYF3fy0HYnQlsCOH9us+AARkm78sdjQY18Y1R9rRzdINGlLuDoNW24p0
0D/1rVTYf3rGmt/hAnEo+3SLskjdxIhcuUMMoVZ7F686Ylmjtx2fpTqasSzeUO7q
o+7GI6p+vA2eT9DBGLWqC8SSlY64ZjeJN9x7yxYxQaGEysEN5kvX63c3q5sHeCoZ
Tp2Lprbll/VfVj2IiG8OLqsNx6RvIddXU298O6CE09p/a6ASoCVtT/GcBPOlNuI/
eNfOp7DwdqZOmqD9brv7YNHee3FFJrl1Hpk1D8Vytr4pKWT/87FxJHzLmqGWIN4P
s0EcXWkc+NiuSzdoGnjePdssRvjwQUK11YZwBbrFMQ7F897sHo4Kh/O7FyCLrY03
NqJPuvedY5RwuGCyULWcaJiwfkjoONx/Gz2lGed/8cBju6RBzuArOH2N/Pr96zYC
pU5jhrzqcIcDA2kxI6HWo/TxFSm+aG1HMqtEzVYivD/OebRxYhSyUyqQE6YCfxxM
FOsES+zlnAIqy7eA/ZInFqj/oDM29PnAt3x7LDbBp4p3P0iljCKYLCE9T+Z2lUH4
e/Cj/W93rgC7tIvbXUBCYeZ599lLrCJMgt/hOEGjQkL7WXyELPcOHoKQY2cEGTIo
1cR+Ibukn3ktYcYRBNoTprOxPYUnsnCOmg9uDLRnm1t5E5n7LqJH6qfPyEIsYTlY
YBvIYvxZ6lB7UxNgohYCV8gyFIEHUfJi5tx2s16GIxqOVFhJYYos5iADaXRE1o7+
CUQeQDDqJF09jCTL6tRHAmXvBhLTHOEjAFt0LBaphp3q2cZhMhATOXF6dD7YQNJ3
5qHAcUTdqGlQI/0aaUuH5QXMOG1uRKlEKFyfwVIqcGsFYqrWPB+lnLZ7XSdM+9rK
pq0DxZ/Qm1WUQObxBSt4JLWjdwJNrbV9xAHTopS9X0lvbsVpRGlzqr6PiPorBBBk
qXpZGb3KHWcVRn4fncD2eFdxB8PuHTApqfUgGPd5bePegAIRrIkw48M2F8410oL0
DyiWdWVl+RmqsELb4HFGOy4KQi2KyZp1vzj4/v/7EvDi0FrsYk2bLPp2wEHDAkkB
rQghvuYqjhZ6TwEY4ft2aLow1FE2Ui1+JGLYsOf+Rv5KPvaukWHv2dVSfl3Wgn8N
j/dualw8aBmYHms66jSdUA+1KGHeXyiEstEfuh/hCiAnx3gXDeGJM8XkwPSq6Fqj
QGzgXEQOJMIFSkKlkEAtilLEd7uBX2I81l1legeE9S7e/f+7iXHqmbO78XuBxZ79
P+ZHkPXIqUO9FEdGtRIGaHoi4Zf2fWa4SGYJZyxrDTf0w0kRbkuXvSypJAeTqbEg
yccMf7yl3wWAIXRpCiys5lS9vPcDlU/HgJ8cZzIEMh4+U57a6wGj0WwJp/rTHvxT
ah8+x2sxM4dqEXH68dOqso0PmRP9DCzHyy5zO9vDqYnR6TR0m0QWC5ktIditABE2
dGiwRPXoIfrUbiJ1JYEcdn/m88WLO2hcvP8ecft57cfZ0MBJWbuoKHqOMHahQkt4
W/mrUGOnaDVug3I73TFseHgT6JBxEtrtpIFHMzO+cNZPXMrjDnS5xL/FIz4HT3Z7
F+3lcHu4hE4eYhjW03gATFRhkG4WOucxXqEdDLHGCSIBC6ZR9FwHUjyoqj4iYb4T
cBCJqs+Cu232+STL16I3FZ5GpFnJFS7hUYzrXCTPy3XO9GOPeU/ql55sQKQaZHTJ
rC9vvgPoP5zDRXe9XnGy0KTLLCxpEADYTXe37z7ohkb/lfe8/XRK4+tnUUv8PCO8
G7tiHJKKD87Rqa+iSThB+VrqS3IzPey04c/M3sa/cYmSTXWFJrDYBbUIltiTY+zp
LTGwONDJO2SveXizagaF/vyZji6cA0MCm81ZOJz8TBQN+MZLI9SVTEos0D69JjeQ
0sZ9zY8eITqQWE53GPjD2lvZX2svoBKa7ewm3OA8aM26UTl3OYIUqK1KDnAydTlg
VXDAXqmcsMCkOhTVoNIiTgbnhMIUUtO5E/5YKGKj0y9YM0gj1clSFmyiZn/ju30D
U++kHZ1EVJZwv9buJ+lC9e2L77MUYvJNU/cPEVpQ7ZOiD3uZblcfl74iS1bd1tNF
XSOXgxhr6U+GNUx5zEYP+EJKDXrMNScXG90aXEol3yn4zQG6kQTW3wBV4QDiOivp
leEjzI9on9+TiCqbJFh8EQb7Z/wil26Wy0L93iX70t+zrkwvzNKC6tAg13R6n3Rv
M0vNtxoy8F/+ow4zMexYcnAMy5WhXWRSYbE7Tq9LwSiqCI+ioDMPVMRUqklag0Cy
acZ77MobhqhXN1b6940V6vTwnwS86fzHqfmGeWBjLWGYq0aZV1p13LlAwohTWrpd
gn7EU9xAqxFjMBwvrisMW90Ie439bsRTbjww/zV5qAyvEx5Q8UwecWBzXdNZ1SKv
irKrVORcZcsAjNd8LNZJWneE8wd0lbwQc9jKJrPA3fD/bOEdIHibB/9mk+r4Yu0n
iG3Y2Jg5n/jR0VpO84k8ufVGTkY1SOa3Kt3/o5OfHQ7niEiWTL4Mv/gvDD5GnSTv
AHvOUIMDnSpHEeSulLfK3Ts/yZBFI9695/7Av3HPA8HBBfwnNAZ7FROMuMa6qRjV
L/UJvJVSfdktPMeCESMstc/g6SjbSlj1U+eh2XOpbsRoy7QCTJH6mLkR1BTGw3QJ
+IZiMUSK7gNjPS3s25LfDS9cZ23Qq0DJtPc+dFtCuDdYFPs78G/4wkUOy7pckdwp
O6pkCIr341hLqP4mvdyXHvtt9Nngh2npw8tbnksrQg12C/EyBrYxe3dLhTEfC+3j
NG2r2/ltyEz/mIXqjbx3Jym20RYkiKpYi3R9Na4oYUdEJr4+nra7Z1KsngxBzvsR
mTir0nzzrD9AFQk91rJUNbUWmqm+2oYAuO8L+9OPoQSCx/l+BCD4iP67ZuoH3yko
7arO5HSk9QJ5Um5J1CPyIKZe5hvyslwbWgFx+NKKEUluXCAqNC0qdH/PUBKKCN1P
J0SZQ0iQEIPFsh7vECgt3b8888Qrbi0rol6yDfflAJwnVsiI9XftSOGtNGJ5jzk1
UdMTWsSuLwVcMTBg22413VIV+kdsd90HpnZqz2M5FwsRTW8blPx7PGz+SjwpqNDD
2IisWbqmKlH6F5Qa2ce/gUibENdq0A840UzefrIbF2VDHWAUm3Pt1Ckxn7nNMTdd
Oav1T9/oOL9vESH+ebvvqLZdRjOAwvqqbZ6JGvm5izJniCn0y8Z0GdNNno5JIDtY
jOMSLD0NfuWeFhIEKcMAaTYxgP5oaoueNoIniuPmtbLJmy+elbEWA9xlNa3lIZ7n
R2ouCcaIfV5U5wFsDkAAYtJKmqF4hpm6C39BfIIjPWn8wKl58QVFz9MbL65k7GyJ
rV3kDh2QkcdZHXDIral9t+kQI9xAM75EA1mxx0xh605nYNLSalIqzDFpX2407MB2
SrzwswgjVMNtmTr4v8ZGkzOzHs/ffZiim8kiQKvPHdXM7r+aHgSfqyddUjhnNvAI
i2k6V5C9QZGdm0xRci6hQqoW4Jkgwp9Ky2JLqlXNcLryDs99S2nZczA39olhjLKN
SLugNWPDRX5Py/Op2rbOs1NRWSz11kQIsBe6jvhwZTSqbPzjQGgtWBGsYqTdPsMv
lnnKAbBP0SKBn56AujXVAizE+HIae9UZKRpKujlHJoRRjTdxOoq1eOpF7ptyLBwW
EqwPxiZ/bLOhL1kwR+dFw8qzknae49bqAOprJsZSvKuyvb6Pw2pm1KFL7BBuee9Y
G+Xel9zjhzf/l0BXo0+TJMqRFOe1xY1GP+1wtVNcRDMkuo/aWtJYNR4NuGHUbrcm
LMGgkDKfrK5FzBvWZiC6KN11Dyx38Cc1MuinXHYsIuKOU1Kfjd17NcxlBQka1JXR
TWVlgSk5V5/2U2g+FsduFOJaOYxpNAlvi2G1iFtAYAME2S1+e6zTzWz9gVEzClZo
SECFQyeZ30purerwAily9ArZLDcdGwUT9tQ63KAD6j0M/7EhFBGi9esDdgN66Vr+
TDNb423oR7sVf9KHVkjbymgcSxKIEFwY1uWAFui2St7ck5FRQU9XW/S1z+wDRQN+
XBdjNl+ePDwrrFRAMOtd0i83peHdEpoen2yo7LhGsjT+nSwh27l4HCVYHEyCq2bW
CRoSa7Cd8QtaKr7V928QyGO2PXTDjbdZqo2tI9XTl0ZGPKVqTbJdztR0anqNjGxD
b3D9PogqTbJOtyJSGM/8ji8tEFBbBO3Y9ywanb+kC76PKIA2i/fTgqn9ECKVO42i
6OS9pW5srVoXXmzcubMrdCKSlV/amJVa4JU0Eee+xPoRlkKixD4Mib0/dgQuDF73
KMO1eX5Ym9h4nlcjHJlUjzsfUCXZytOdsnPalXQe/X7Ahe83AwsUE4B9QWTUke6y
O/BUqL57y5GM5TvUak11QalrtX894AuGB4D2ca0r24nRTbzKHGY4J4jaxd7zHOhE
WG8a9SaJbieR7Uvv32KNpUfXqNxTtcf6vbg782bs1rJGoZPj/d5d6Nlz9L78W5la
3hjk1mutiH0YLcj6ex9FXo2gPpUDY0y8UQlqxmvoiJdtv9qyBduUib07s8yFC0hG
3WrsGlvbKU9D+6Ok7juI2ESAU1ZAPeAEl7+YWsjZ8v8zN+q2gPs2abK/izvr2Ys7
KdGLgYK8t2wj9/6ECifPjOznNzK0lTAy1M8+jvGo1Go+kAt/CZdJILjCTFBmt3pf
d52N4V0yLBtULkEopKe0BslmwcNiW6uW4J36jDqYm6jmyh1tX4abED3IZj836OxJ
USl/N5mxENs2QBFWZlFYLBdS0+b9JmJrNwh8VZk07wjkKrQxJlUOCAPHXG61i/k+
FCUkNi4SSGc3KL+rnRCdhttMmsViYXoX9v5LiAX6MOMiVRXqMgnbWaXNOSbomqe6
XsS1L9sKgx+IDGupHGdjPZ7/ZDo/OHDRVN/ShSY52wlF1/HhnQC8Ce1XBNl6yEaP
Q6fdXlGWZjfXhxewadPY6cIkv/k3Zq3un13ZiYuheIpWJZHPUXkTxKkzFnbPrzWt
GWtFD6GEyVQv6oH6XZ11Ik6JArPXeGvbhK5E/YL27tiHO6j0C4x/NgR0RhKhyCoE
86drv023Lbn49TfBTHYb+B/WrqgXcF7Ugj9Jbl8f5C81/ZGUNBOqvCpmKSsqo78F
H8xjfXs03Ho6jutHazmUh2KZY0SqpDBupSM8UvYytIgM99mvMIbq5b9Trk4beRvb
b9uHa9uBf8na/QRVZBweNgUWVnWoLu3AykC9b1UqBAq39m/omWv20pd0cPvmCZ7I
QqmF2hphkFie6LYMZsPbEf2cx6lU0x2n4SPWCU2vjuLcbT1DFeP/k3ANg5jJNvAg
NjRbWVWtnKKDDA93kKWoOFeYgeUT9lYdPBbVvC79wTr5lWrJXH56iiZ4AYuOl/sr
wfqkVIeuzf10cS6LIcZ7eevK0GWA76pm7mnRQ7PZrhqYH/Px+p0egFaGeqTS4o3Q
YN1l4cnorLNy5XbOQDwahGQe8IE8v1CX14H+o804VomfW5s5NjUw3df31RvlKuGR
zySKWBRvvdyCfvy8HRqMIR+JA/tdl2Rr022E1nnNKQLXIJtOdyqafQ06UWmWx4BU
Uioi77t9w1jP5+LfHMfB2ssYWFOtPJUQGlBdC/Bh843Qw92C3TYoW57kZpuHeei0
fkII8UmdwPFFK2dvTcmf+4GzKH/UoH5OHgQvucfNO6Kig7FlOxuE1GH0rGfr2OPl
IXHmrmAct2KfheLhnx30tlztXLCWQ0hsxpvFcMwSXZyFUwEkskMB1PLIdcQsaD/E
7auVELexTChrSj6F/8ytsCjgPvK7kw3HxVX6Xng9qZT/ilcxIigaQfu5Srsc/C6v
t6s5kNKyNCmXFzp+51FkEgbHJUsgojkTSov1FBnWl3jqIvYFyRUaKFitGRfjULn0
HSAxA0qIinhQtrRggvG7Z2LmzI2VAkG5i0D8H0UM4NAb4qhYFBtOVVDAG58/J91T
xImd7+AbidmNawWVWTjsHR6e6oYgyUxPci4xqjgaumqy3w1zWdDFMGfw+XANs3wm
qevlK8NScgbo8qqi60nfQlSoNvosjoPsb1Z7JI8gtcnIkUDpyC1gHw7hcfova0Bq
6CEoiOowOIHzy5t54pkd5D3V9cITaO+z5gbzfOTQMm+WElEfKpZG+XNQS/+w4q1G
/JmLrRUm9wDuI2QocvJ7i2HxiRbjhg7Jen95sUcL4DhS+aVNWtoJZ50ibPz/r81+
OBv5yeiwnqk4vrHgUispiny3JYdJWRK1wV6JRKiCoeP8/EiTfpNGfMCCo8Usy6yE
4J+5EFO4Arv0fc1voTsYKgERX8wbz9l4VPUL7MQPwQXUprrLUcR/KQAW90Xg4WhW
mXjRc9QSb9WlWzyrAVSCatfreTtZOUGGi1InOtFqweMuDnBsp8JrqFIZTvW/Ulbw
Y5mBH90m403Ol3BFH9PaqobcZGgr7p1EMEDfuv06RqN9Tv84kESjdm5RGUljuUtw
WAOXMYyn3v5nyfcXn26Yz9jTu+F2odLtgtShYG/cWElh8jZm1QhD/aCmIJRqTDia
bUXGA/RjnpAJ2w442gkOnSGDhQMMhiukcY36z+iQcZG56GW/p2Cs9HzpwQxZtgkK
2MRlrkQ/fv8NRFVbGeFVUiMSv44oHVscZZVMdxeHXVnHSxUmJs9acKRbrhSJzqDu
BVbe/i2xYjBokiHDZFOSsyCAO1e/cFyEkIJX3xbN6O1aMq4vXg8pIhxjM6ITXzLg
Rt3G2o+ejgfCxbscrhTF/l89HdySxSX4PSf5xHZhPVgB2QVCavXtMWMxAzL3EV4p
YTO1wlrHe4N9iskVuENlOpmq31z9SSinsTDg52hEdUXJEJPix6ypIKwdimXTUeIJ
NnsXS/r0MEhL3yMXIA4FJ4IWXY/c2149DPurr3WoJPyeL0F7jhK7EmKjGtPfUOoZ
oeb7HslAOtK/zW+i+w5aNJVA1aLKm9SLnZfrlWyZxeucXSBhPbZsuPDI8uo1JKUg
CKWqR9X6d3NyvUtOiRmAI3Xp95ofzfaNUh551FNAic7nEQKH9aaAyodRdW+VeTGi
0Og7M5I1iaGjNuMz5512EPMu73gMUlmcBnNUN2uZDlgCyL4ECsLOkl5tup6v6RAL
BxVQTm4SaeVt4JXQkiZAGVrWNUriQfXjA7wvNCRHYomLCUMSV6MSvjox8EkNAJxz
TvKXMdP1JNzFXwbofQq4dAPCF1a6npthBZX3ajaVG6uZIlx+HsAeLF1YXyHRFztj
puuswAM4PFNOgEnJB6l2HsuXpWB1n4mD41gaf1rcbU8mxHZmEFuXx3HgiM/OM3as
HNbNOxtXtDzIJ/dr6ITBS0aiLopyf6Lbe8677DRfBb+yzoDFOnOZKjo4vO7o0q9H
PT+aCLByy5+cRAE4WRbMNfBMt4IUyFLgkLwsJ39G8KZSh7VAcbVfy+8S6pRBlnqm
EemXyQhpIi5vD+bT0mpjKZIxSZE/aAkvVvYWXByls/nY3zF/rOHa2x86L4iLDrip
wOM5+iJfdztRN4pFeB4ybzYvosWJ1RRLXwAyJSSrNjLeLulCEFj2kHp/Wpm9lr1F
Nl7wijbtapIesy1gFMoGC3SHInYa06chTB9TEHfhFbttWIHTxCw2g1ek6tv+V2Ju
b1eva7GoxZCiobygOEyWZJUapWAAuF60RALWTM4BrWhRFKvRFILtS76JEDoKhlZ8
i2GhpNxpK4QU/aWdzo122F/gpJ15Zyo8iNxIloKcRtSCZa6Xcct6wCbKDxynaFiU
Wis12jcJdBr/ChYL0L9xNkqL+7ZvZrzAOXvDyp4iIwa14VuHpDHitSYYRBznsEEm
/W1J+adeftMBEGAhuEUWUwnIH7ciggcePXi/EnqOE9NWBYvbPWU43eLytB8pHp/0
G2iNhHevGudIlqr1CKCuB/iJdmAL/r022NaaPIAtcuEdxBIMmZZxe1vBq8rI1woO
E/D0I7B91Tw2rDEvxJBUr2qum8zvXLR0XDemb9U5VvFflOpYGKKk6j8v7sOGSPsu
CyI2HrG6QTEZpFUPkHHQ9afAdlxj1sJHr8196eULPe2mrphNiXkl4iLUfavIMElz
IuwQW0qrH6G+on2Qvq08proWopJk58Kxv8iCdkwkOk8MI50EcA0ThL2MaYnMe2ly
YvgIujx6g/IQE6ADFOxoD13tOFfE1ZQWmCEmysAVWpoFbfmQxdKgimiLArjSRxKD
D+42u7K2BAqQyRAv+tOYMXkxqL3FnyG30tAZX9v8dQnAg43xZ23j053OSBSux2cH
mnz0CExbxNNGOhNvwieDdGB9u31vW2xNa+UHtnO8Ki+rVz5ZJspqQ13JQM3oBlNp
q+8QL6kOLcNGRDoBxWjzh1/OEmijbp7J2+dNPBnse66YzEqManqWX+3/fN9bmy7l
TDe2vnuwWBNHaxEHdCHt1ol96qJI0W2szehq5CPBt61s4ytAuz6BITirQH0CqXjE
SXjRRArK0oCbTNWiqtWgGOA3qD6vVb51zO8RRFX3N36ubDgOCVPExZkLr9kr5Zyz
qiGowXbr3Pfzn7SgUAUuxMhrmlgrvgCzvActiosdf6Tb6C+MGcVjoPx5+I47jXn4
Pbrb86SF+z5WT9JvqXV8+hB60w/Fu1UWKMPq3rsipyNOFNxVVCMuB4unRNyPJ5+c
g9hyR5TFJ11Tw1CMBIKfZ5kPnvu/TZSii03wn+MmmB6dSjydrmL7ZPVvyfH2Q8pk
7jTEiYuz/N9Ghd4+3+dVOH0tDyFrPDDp3iBUp7mxPswP+7cTV+WVWvRaXofdDkLL
696ciDI8EO9ehsNTVWAqUzbXVsfw450/7/pVV3NilORu9KSI9gAaUoEaU3Zf+VP2
t6DxiOzb8C0EwMKFGrQ75bZgeIABbUNimHQvCxb6dO0hvBdwKx6UPGTbwCwC3Gr7
UX9O6yY17Mk907kzL1L/hnc+Zq8yLi7V3IMGESm2Ud9TCz7WuQkj1cLTFgbJTXyJ
49r2h2Ln5JLBngBsC8DTFX5lWK4FPSd6Gb1X5slbIysroADmL42uTH81G2iQv06F
e9boGNHdkVpSlPnn2s9dA9g0f3/p/Wm0O4QbJCRL9UKCC4D9eQDkqTts7s46CFdV
84I9K7p3kK7SpfmiNfHcl6Wbq6VXUcOoQO8phDzOZCek0CwFlmMXpYrHI21JX7gQ
4276d+aMj/6+54p9MGmPQcoOKL73NKsGMtgEN4NuYICtSTgaAkyiiPSSif/AtAYT
PKR6AIEWXjYiyELKmg40AC4WApqH+f3SVZ1ag7zfK+An2dullbtxHa+mPP/Xi/+s
Zly7KmUpzu9F+KoM+Bb8FX2s5Ac7R9WY590KQ9rYpK93iYrPiNR/fG1eQKsdqjkw
lf7wF1bbsB6kr1V1rg2vOGu2RC3SnzIVm77uO13j1u0F6q9sITlyT4aynBahWHvQ
ve+IUQSL3mgJwca2rwQOit2Z4e++Z8OjqaVfEmQ8wbkkHI6PPqrN8UXMTCcg5+cM
i2pza8c8ZY+yQMJn9ClOWoTA4HXSh5BWPxHC+/Z8PRbDC+0Dk8Cf3vnl6gF9ZKr0
8g8BSQSsWrTr4FWx+o/+0qpfGGgsBQ+OlXS77XN+ZTV3rBzgQ0Lxh83/VaQdnMTA
X761z0or5jTUI/h2iNEMFo42eL5Cz5RPEOZS0YQgDcCL09O70xuQurqky6jOLjY5
UP2xduwsgactUgfOdbV/EiAwAQWlIgqL67fTKKQVpM76DMXzlsCP9ILDBCQKgRB0
i7E2DjtX7vKgkuPcUw4P5s+8wQaLfhdv5ByLlYaTKIe57KTbBML7mh+Q3juKhwSx
9N+fHCJffc+HyO8tz9/EzCDgts5kpfs9gPBURCzCrz9vWU7c2O+NvGVZ9dtZb9wJ
1aLOPwkqMYjumLa0ohN9UAJMbGsQvYvkRg3sejLwNilVoD4k2CJqld8c0CrJk7UE
rLXdJqeqDBjUv3vvrp6k3duyoHaw+JCNlriTdf760z0M3sCXwW5BKxFXwQzX6sRB
fdGg4cmJXiQDzftTOkPxEZ/PV8FOjLoLtuZVZN1AODgamUlmo3xMyZaVDCgcNkqy
Eo0/U5zcJpRWDlKUGhw40uJvqttXqt0cJTu+f7LdRVZhx+CnrpT3rg21JnPAPxLR
rDx8i39nFjE5y5eEpoc0DKUqHc45EKN4dXw8VjcspGAzAvsqW2nnAEXNfipMkj0T
mb2QtCmFg2DAy2G/BohzUcrsJ5NbywVNyMnUK4DUj0fgN/t5CbeQWKyHr9CO3M++
hZ3Vg4jZWlFe89WOXAonXRqYk2IcHxnCltcJHoHwBf+0wz149WQBdD8pqUprh0vG
hh6vPOJvAlciO57vWNeqIcl0zFAinCaj0QrJz4yoarxnyYxTn7MHX7ihLxIpZXAz
AhW5E5eZiPJYPIjh9f8CGm+O3fCDq1Wi/JvjO1aS2B5fgZUEN0gM6IynfHFBOaca
ui2kucDHMU+o6638Y1f12a2FoNbhkxtmevIoRp2fzN7kew9rHEy1WdOYBP1e9G/j
DJ35n4sguCz3Jm7mXwE6OlfFxDwp7Ta3USkXWF1hSf7HpcArgA7DaeX0dYj0l5jE
XLpSLyJk0avkzxMSdNHAIOVPWzeuxSnuffcZvZWwP1fI330T57qkWSYjskzKkUDG
bs7PuivMPJLWe9F6z0ZW/nCf4/ZhpRFewLLOEs/zjO63SApH/j9zS3US/xfUtyD0
x06ulwDQt+T/85nWeT7y3R06bXFKHlOi3Tb7CCV1bqcNNZHG1e/GOMntAi9QZWfr
IAn4vBJCFhTy4Oi9BE7LdeFirGA6WTH3228qCvz3+4bbB4p5wObBe715NRaE5YQY
/nGdCGlP4O4rQvKu0RRX8mb6OUiEQFuvO5qc8kyqQ2YcAJe7244MhAIG8fadsis0
O1sTAUgzTuWxf2dkVjbjnwUmAcX2DPILYIz+OUw1/iUCfKrkmBaOo9F+XwzjqreT
fuogJK1slPYl8qWJFiVuDl8i0QhRz4SjW80Tt+x+s1SCvYcGQFd6gWclW7S87Sls
3Bb+DpoWojPqmjH58g4xIjdJhH41HWkq/L4lT12Wj4AKD1aR0hudeS8HAohkuZjT
2PEX/Pxah3sGoeaMc4Gwkgqo7ituZoRwOVErr3gq5h9o0T4SC+arYGLzQfw0OQq7
G4yfSZLIrC3ePXpTyLztDO0fa++3yfHIWaKnHSQ7Gblcn5ggmXdOLNbDE75WiJiX
KrF09rj/QEKCE8ORzlAxAt9hl9G2MYATR6RJ8tRnK7a7d0dEI437EXUQac5Xm3FO
xT/FgmMPZUIBHvT2zfIGQTRsvPfQrWl6lXl7LcrHa+WEEQUCeXWmHc2MAZIWdipU
iwqviAwNZjtuJpg8ihPBMHPZmRBqdCN1qU7+fVJ0gUnJ3twbm+4uyFJDFN1cYTAC
/jmfbd7fPmjhb6GdE4BHl8v3roNFwhmGyAajPXeQl6BL+p6mVoAgmHQsFddjO7Zx
km8Bx0YIaX34Or/IqEWcjBDRxumbGXzmqyzhFph28FoCLjKtikH4J6566bdeNkvQ
XgXgl3tAyS9Tkdn7X7js6tCaX2em7o2BkwS0Yp/Eaqrip+vD+OAPArJ9+P65AaOu
w3ItaupggvWIM7wG71P/OFOx1WrYVbfN+oy4eyO6g+FtiuNs6B7id5EoQMA9UwSq
qhZxs70mAbmtDZjanfqEUo8YeeJrwyyMugBYwGOzSAMleDa2TP7ytlTwRfdFvEBp
ureZUNB05NmxgX2b/REnZkejQsFbsciGPdd0TqepIwR72XT8eNui7C7ErYBsmZmA
o7/uHwmG2mxQ7XZsvZBpgDVVLag0DCov2c2WtaQT0lkRLk7XAJrJ0+ZobMkIl+qs
XItN40XEX+U3cMKe38Xw2e1qFpB9SQmdZV9fhgfNGGS55KApEp20E2lMsFBa9NLF
B7LfMDOstaR/UkjgehUeJsgG85yCf04qdfAqJnr27HGbTL7RCr4OZOxW5YQlgUBE
J5lX65WpqEXaLwZmSC9QRHu/G8m/ZWm84L19SiNvg8GnB3wHQygKgICL9d5mekSM
YpFhQS5bXrUvyHqP5bBUDLZxgY4NqTYtSjlpcLhz34EyX+nMByzTVcKYhWSduIQX
nKywX5wTqFpUSqKAqZgUFhhtuJqdSCgrLyPW9PDLrIZOw1r60oZdFrV7vOkSjOIc
p6LIqZvwQsK2b9GOpjmn4zSMT4GMa30Di017iAHDkmgMCIkiLH/7ZjBhPnoJyF5E
DTXwoejo2/pvB/XZcgvyn6Lu6AiGlOPEPJBYpMhjQ/ZQxxj9yr1UCchiJGw2Gmto
wJgZJrIQjgfnw6S/ZLcqX5Aa+kGNEkLbnvINPC4I1i550FscF+cdwk7USDn8dNiy
1k/mQrNVl45rdhmVmRu57ODuJ0Vn0fhQQTi4Ah8fhUNOJ0hl6EX6KJtGyl8rmzGp
zjmAHj4rNWwX4jYY/Adpk4TVTXsRCE6iMT0fb+X1tIAYU5dj18D7j34agrCiMGrT
Lb9ypqF16sd9odo4E+JPO8bZ1Q6cu92nXTJoOXRLF4VMWR7VM9zIuDfJd7/2qa5O
FoBxJ4x6qjDA/82sj9812tC7RtWMJkturRfjHpiBJP0lBATqn9eNE8gVxs46WO36
fdtL7BQAHw5+JTdHCUK8bhfF63aNav9DITEjKZ1epHGknT3vEr2y+B9c7cBWcD/h
P4PYJNgjfhkGiQkbSIgjtOA2ox47bv1GrxYY1CRQ/vpXu0uYRLOcjnkHoANHi3Pg
qtWplCxG6xCjdYX6VwDucQ0yVlHQVloB5uBjWENwKnETO1DAEVvM7vTzd/aHovwZ
inBDelzkMiKdKu48xu7LOf7hcxAPYta8t84Kyi+jN+6R2fega+dFkN4RkN2eOl76
uAPEta3NJIl0sE8ymbAFylEBuYvfHsgdBmpyyuVycOARg0feZRcIM5RojapYiKFv
dxEBoIzwK3zD0HzQ5Vv1lF6nNyhIdP28KJFWfmMn6a7akh92utZjvMn5HzPKGWrS
EoxfiBLuo4gYfZISgMCcs8dZIXiv8BCoMjrJzQagfLk/nhjIUb/N28k0gtsaqXdq
B2xK1py+uxznBnlnIU2pWPu0LQbiOE6BiIO9szywBgKZXFOo4h+3m6NfGFXO1Mgj
X34aVxU20hMkofBj8fGw8bGLeixAWMsl+mLijWJ3wEEa9HgQ0mkGPSDKb0okEI8o
L7bUAftKZUw6+3jwSBtKfmQNCyWg7KJDqjSLWqppq14yWy9BAQtJgKnTUg2XglIO
ZyDEzsMyZUzFUA6STW4LTKAQAtdpVszboeHNBsDvgct7arK5xU3kxtLg4Llro36n
TCcMLlG/m9dkkVt1Sxojps5Ze0oOrr8x8HusY975InsQxs5RpwTzaktBzRhEGaoq
HtCC6YouY6yrrca60OJ1nCyQu0YudaIN5fogl5C2gfOGzvs71iZNAzscPu7kt0b6
aH+bs0AheO80JLgdFHtuAA/BNhcVlaPU6vgIh1TRhVTEQXOY7I1C6k3ZPXehSm2Z
CU/DtCuP+Xnx/WXxF8tNLrPdOVlEHpGsv0L79BenMa8x3eK2DUBOZpzJ0XTYxoBT
pZI2A0RGNGuq5w6MkZ7uZE4uwNBDjGoDq0tpT3zfhHN4dpqpc8NDAKhjbOhP9uSK
+dgoqIEa9svUno+150fkkCPKQs+0Rb8WRQrt+QIIMikKYAaX8WgRhBhAgyEYBAZV
ks4YlkM0wuiW+3J0Ougrgj1yZiKnn/UIOX8JpySvzq7ZOnjCPkYI1KjdIYSUYv8F
6Xcd6mgfPFWq3gfrOgchUrGmklqfsQAkvngBNXEaz8iP+wT/HX7HCTW+eg+L7gEM
c2Ij+I0jT06XQT0iCQ4213VSb8w0ZFfTcZLAwJ4mHRDDz/8WAdu8JC+04R7AIrfI
LIL0j7IHgb3iNJVfmA2nAAYLyntXmDFHfl9m9EZIykn1x9MoLqdHniBeDUqfYNyy
awJY9iGiU40Ysf/IuLPP4vVRPxnKEqSEn8dhpblNRuNafQ8V3asqA/7WFJ5fL+hw
hQsMDujpznZ8nbikzVSsMdDNN2EC8avupseDWNff+7Wb8xCwJTOL95GASFCDSD91
KWfZ7KUGGwUVC9jWtMeSkxs4TdLmqANqTH+8LVEdJVDUYaDG2rn57Mp8IMiHWsIu
5jgDbwaoH10pBmt69UWP1HdxcH0vStXWeg5CyjtmfN/VA/g2ExHLiFvR6P43rwtr
YH0VWzMVwKZrvuYES4zYVdnLbOBmF/88jpcb5tSANrs8f6YEKRhMXuOTsx/Q62Q8
Iwo3wFhiJFgPRZveDYIo455ePrb1YGPNs7mMBLuIcvCIlaiwixXJ4xoG8GqBI1xU
qlruTxrNsrcN9hv9e+DQIDIKo+a0BmQILDP89fFxutwqseQ/4sDg/5GgRhwCocIw
oEixKy4aFqD0JUxsOkVsqEg97CKWjowL02Kh/ieRO3l/aa7qjVAUinAHnxVoTFDo
+ktzFrnkS0FlE7Nlcf2aB66YYf+SSvXBORrC9O6WIJ2gQAstznPR0xuaMz2wf41Q
aNVW/lL8nkuLal8P0xR2SrZ+fyIY+LJ2wGGuPQPU9yCwNV3XnkPjx7CjzmYH5d98
wZxV49uSxrsa4wWWgclTUTu/yyNGPMV02uewM1MVUPCTVKYbaWuffRRrfYwP1Trc
W8c9ftYB4KDomzm8CCAUx224ZWr8fH0RbLxjlJ0IQljeRz5tmhpqiBkbMGMVanO8
NeyrvJ5hbN937Wlq/xZn6TYFbACHSx0dAh5/KveYRMkb8Ckz4fdKEdKGQWgn4+Zx
vQe9Y+NYEA7Rg1u6b+bnOgHVedObqN5EFoMARaxrUNzJ/I3GSjrFy8mZ+s7fIewT
0c5gHPGBOP5KX+/7Haalc0dvTunfR3AurBP48pGimvquwK1CZgPsau4YWGUjES7B
OEwwIQsgyiSpRCZXkle53gRroJnj2AwD71nsf0BL971a6fVl6vP6PmUkR8DXVQX7
6l/Y7IlWkQCUurjanuSa7fHHWNWOGztmdzawEe2zRRf6LM9XL/kB+ScykV6IxT2o
+HvVfvzD2LpDxtTluS6FNmfw6FRp8QxTKD/eNfy2RWN2hmSiQscYXslAm78sKKCz
esMyXtJkgag65iDb13PePUKRU99JRc96hP5H66G9nqdh/tz6Ypwtn7GOf46Oz/NC
afFlf9hNH1j38DfBMunHEavdKp+5sLudqLtMbcLBhXjXN0D6SIpGX6vtPwq8mV6y
mtEnV43whi4wQH7IN9sAp+pFVGBeFgdN0p+rIGPhUpqamlK77SEM7gg+xrThYuEL
nWYM8gUYDzt/SeA6CQNUSyL97tisjU2d2tspjJLJNVK1zCV667wn/2l69qBQNUa4
PbPoiJniMPWxjl8w3vt5CbNhNgDCMioylBoC+zKXM2HYemoO54Q8psbcBESxqf0J
ebg08akziyMjbD6TZImphds1pJYOKvOhUirYsSghLecykt8C+2dRp3PNiDqUiGO0
pHKloKvvyCYD4h0UsAKIhEzaQuTnP6czw2ZnDOdmVnPZrnPPk8fnhX46YJBGsT6F
J1yzBD9bvABn7sai0W/JPpoIJqYMkLaUvd57560eNIlhjupTY29a1k7YLATOj0Qh
r2PiBe3QupkFI6MiJkemXEXaD/KUSvR/rydMcxGPQlsg2/ZFw5rLz+JrGQA6aNWa
9rpFCzKapVPzX8tdrKuKHcvMPELqHwYGns+29T60M8JjzBur7YCrbwbVc9LxSy+j
epu62m8EKPQVtCFnNL1FlLmAxMG+DmWOy/qNKdUXdDrlC3cqIdDReV6vAr+EcpY5
qeKTwb7QDQbLt/ir68emA+yTfXF8JMvkdx9N0nf8Saup1WuDpGBDVaj1FGE8k+yd
qV3uR2Y598HrvEX0QBJD7cEInsDuTTpBXDK7KV9Au0wtjoSBa56zyWaRu/Vg7yTq
g9wK+9YutgLaIzv+hNa+6BeLfMeheEq28naHFkppc93bhMs+pXDMY4nHd4MYKete
IqFmP8kVjuEp+lNyCln4qB8AYZR/T3uYNfnApp6WQ6bm+ebcDrn7UnOVLvMSuMzE
lX/iT3eVo7zBKXZ0ENYXucF8C0OPDGlwacVB5OzlcfnmcHQtLsfO3MlhVAy95PMy
R4r2LTZkjQFcrTATRdLSb2lqnyI2cUqwtEUpwWoxz/pOszsIacblZoskIFuzGUuc
6G5sExr92hkFhUMhKhIaEGV2x/4+M9DnqzV1ZifrqPmfNRB6yevNkt8LPqcpIeLO
x3sj4yRAoJm4uLWg+4xEb9DvihFP0NQ2bcD778xpijRzst36DWDS6D95Mx2Mv2dM
ICm0bO59yMzZxjXsN8SDi2VPb3MFuqjgEjlIaYB6G85tLsQ/AkyAl2z0JSqtzKZh
2fTpV78WDpFf89XKrm8+lqv3v7t3Sw8fwIosKYdY+vhdtQ45OngMRTbTzLRRpbGg
t82plHaZ8f/07efVXmfjt7/Bwrwg/bBr3voKLBUm7xXSwQGermn63vGA4dWjqOUi
BjC77m7N8Uuf0uojzMYX/EiZVqsOdLnLms29940OfoIZ5Eo3gHAlYaxNhppEPJRU
DWJ8ww71MazTI/zMdFs1TkdvzVAAqB/coqB3iUjPna0AV2KCvndY7+rdgCWcKoYr
5vNtJ3zN67uBjC7GpdKvU8nYYQeHBBg2vHHllwQENblxtcBUfOmLcAZ4MeT/Quaz
0kwrwbWJDo0sm+6zezQnBUrouUj3NzaA1wVsYmFGmJfzUs3E0zM37UGVXuTwlLrr
+MNOqrmij1j1soK/rzDgHLlU7aASQtAyboWe9xlwaNJPw2YgL7/aAE8tcEx45mBt
LWUDtFgSbh1kI7hW5ppSSVW44Jl4J65dSsPQVRuxjFWs6xBHCERcqrZHNgzTkF2W
6BwhpMw3XV8DvPQLk/RH3Eu54CD2fORMX//8TtMuVGKteF7xFUVTxrTn95XX8grr
65x3q7LCr3IPuQaGQZIQ5if8XXLyOOpFB7/Uzp0xmsut6vSrLgn231A9wEyug/I1
/A1g/2U4FXNzPVOoSTZHwdpiVlfQWCQYOU1NJIdpo8/dAv7QR4AdQ6semcHxn3vI
TIc2Au2KwdnTBQZwz8wcr0VLwtZlCHlLutkEFmVYRVDu+UoykBjyO6Au3pJgwutE
j2FNdN74uvubxYlT1Vd80BSjJr3BURPouhTkoELHfnfvQflUSRDOTtfEBfucp9wF
eRNjEtLOKbYyJJBQyecC2ieW296eV5mn0PG0K+ukx307G4i5G9bLdxiB7NqRd+Dj
nB3gzA++sqPH9TgW6f5EIsxNYhHwTc6uJVKc8XpCGfxrS6yDsvPi8sR5tmaqBqlM
U5wH525e1dWuI1A/JJHgDkBQ2To3YWAURtFBuw4BEBerGnLXoBaPT4KX42PcyCUf
LY4e2/xp4XygvOjjtQalSv/v3qYfqJjYTfxaI+F4shPOMJlDP7ZxekblBt004R7A
eVk9hhJbmCaIXCMX5DmCllaZEz+jpMWQ14CNeYUaAPtDiE/lAgx1WFGun+pBFyd1
NqVaXE3zAuQM/NdtKhLGHO0C8QOcZKDFPKMAwrh5joreknTHNoxa8n1OsvH0m9Az
ddkVXkkmAmBfj8B/yCuXqdWXcGnjBdxp2A6aiGo05VvF78XCE99xcDdVQnGlQnM2
nocB0ybQ+MAwkNtQilwYzXIlTyp8FUbXTI998RkxNhNHAeLcSaDGFfdZ08AozViN
Qy4GjopcJGdJ+b19eu0SqhDJvy2/o4bKB86zB9vfEo6IOxD0FgrcfjSwskk0p6Kj
MzzKoI6ffQaVe/eI4xRhXL6absb5/p+kjcKIbMdfUMAcsLOyUhYS5/fX0YefWT0y
Qw8jZcJRArufd217GrUHDQz71a8nbB5dHVOHPFzFGo1Ok1Yb9i2v0T7Qu/iQvF6i
Kr94cFxm97fwqQbNznhqzE8T7H2FB9dQT4MDKxrWmeedYcr8LIr0nQNfxgvcHzh5
eP+iGdjGrszEWSDaxiOchYO+8V2S6kt38r2QgbWse2Zp+fWLZI5A9cXUHRk3AiSR
VQZVr6//Ru4WkzI5MuCTlZnZSm9wrsAuQEP9qv9IMC9F3zw4kxA09JVt2Cf+XkN1
dXMtBmUlXJNwGA3uuTQq2QKe8fQEEeF3hWSTRWIqfazLa0NkvOIg8JXTficfJbQ+
0CLFErY8ELiLaAcEwc8v5QUwSaL5YCMyw7Npa/FMTA6oPMVlPiYiezChL/l3bO4v
MLppUcjpYWsg2bgFLn1xptAWsnDzUOTRQFxdP8K+SWklKw6ze6+7QZ6Ui7lajOo+
fLHYrr5zT0RPhYe2EACCZEO/oq1BAx4CqONPJlurIbeg7rvyyKUhSLJnSpMUeH2p
AGokt8+xq0fJr3y5apqwjJGfn0Ze0Lbsco6x2mdz+H8t2MlTJEJUmkuuUi7Z/8ix
R1j3NE+idqDnIWttOgGKt5d6G8XiQjnRPs26rncDmlnqiU9zuDc7gHrNA2BZmSmT
kVR++wmzpGA5IgA0h0bRFoRaA2DBzpmjPJXlWM0giIydH2IAeNJhRVJnV8XYTg1x
1qHyBigcDrIL7+5EQXi6Eei9w/+NZsJ7l9wakW+InmdSEXDYcJJuZAzHKG3bmEaM
+7ktPSDtt2DNqvsEMoS4qIz+DC9FzU7tBbLhbeeldGjVVpOTDP7xTtzBLM3oH8F1
3leD6HhSbEpaohipa73Q2Xh/Er8Aw4oDm1aZi7bul0jeCGBmWUjkRlFLhKBfdvHM
M0XYoGOYb9jTc5mPnMcevAQ6vNT1gNVRcbrFJN/itVA76nowAhpHIRqXv7z8ozAu
/nmuMtC7bHOt7fZsXsmX3r8eCcB36OJ4C1RQyl7q6Un4gkk8pnQUo2cYYX1dDERo
jKgzPZb+PVzyiqCPGkyBxWJNWfhpc0gjBWeXClDaLm+TVJN3xUvp7ZD5ShAI5EC4
Lywy0hZDzso4mB4LMounukmIWfea7JyIT28SivirwwZ/NN8qIGXxdI5rQJPBwpgT
2l8L9qG11Wbr09Lo3XLBM/AEkxglEutCAwSVLBf++JMVkpnIWcS4nc9X0nXOpEoD
IcHfZtDCfV4J/su55imkammtLZUltS/fV+55uAZSFCZx4hbJrNqofCy/qSsY8rHZ
MFyWFl0Ata74DMSmYJdZWkgTGHpYRfZTLT1VYIo3pNlxCnTX2GiRw3SZmiJuJAja
+QYKSYkzMgKRas+Cls1EpE+5Xjl7TWLD9neHppN2jzcR+7f3smypVIx19qEWttKK
AUMsGDJ3bmzx+KgyAKIBKlCIcOqCAS4wmyy3rPC0hbMwwnNrDzGUpYFRHIcPq9pp
vBhy4RoOpK7wCGP1MkOgMgxZaEYieLdRvVpep1vEA5yvx2p5hKMNpfb+TA0Ja5yL
4vg641PHxtfUE/8mdaAG8QfWr/ehtNw+sJieH7F/u5rRMjsEDiWwuOckRH8W+2Ph
skvndssIq0WBkwQ9hkj4xNsaMMO+XSmM1MFGkiWsSkKuyZfX300DKfXL6X/KhQuX
PlrEaXlz/PYnFN7R5wFxQ9kmt1MiiFizvJZLxVijG+20lXxz/h3IdGv2pnkHOgq0
OFG/VDgBj+JSyFRYv1xPv84hPhQqRU+fQeM61DRk7jrGYWvxe4hUi7uozm6lzIxA
PfIsR1NFsJAdqVcqMvw4B2dd/SR7nvSoPa70NpK6JKJWnSTZ4cMh5C6w1lQ8XcgZ
t+d0yQGqddMW8BEq8ADCkYNS4vm6wH96zSe1K3kIsFC8tGProLYRriSmE0jGfo8U
+IziQXdPi949R6XvdUo09XWzty2n21mq3MwtzZUruaSGjuQjMeMfkYBxd/wYxnCv
P4khACQ8A1VocBWs9DpdRmo6J71kOUGq+LQhAmiK1qW1NgPuzpcdYDvYTgy1LPZv
CbpEK10MVVD6UtQu53O/vL9PkJFi+a1CMf3XytoLx3c2gjzTjfCATv+BGA+HFzwO
pj+I8Q02ndpGvCcLS03OAl14ZYJKCE7q8/oLTNq9Wf8zf20iBHc3+S6D9k5GypI8
3SmvqZHf9/whRzKqQQhCR/VAtBpIpAypOxY7mw63jD0hOncP7AsH3ofE6mIyElag
NWa0V4ZrQAaTkRnbkA2br/+RjkXk8QpGccoQfMiutkikJPZW3uRvMBT0RS6U+btR
+dPL/+QgvFgQLPl49ZRts1bCFqluzRqNGZO0AeggBPiKXkuwUSYZJZZEYfV6d3Jv
1uqiOygMo2y0UDMklZlIUBv+6IdKofIovmR8gUQtKzOcK8l2gDP6GHSVRJbr4uE4
EfUp4o3HBMZBLreysr3y57DDMonDKYWXLs2+8hN+t8y11XxNj98AWeqkOa/M2YeA
SJpMd2cSjlmJ9F+BczzOSmXLQQD2cu8fL3rQOSAaOJGfVtU8/0XVm2kIugHyqPHH
rDX/YbvlLJcby9OtMs6SfXHDubpvKr4cwMMY5HUkiDBDT9BMDlT7iSM8kjleKd4G
eEFJMXGZAyVcC9ZkLLLYQ8AdYjuS3yCQ1/5Yasg1s5+0Tq0MCZq1CiOnuA9OyGxY
hPg0NEAe9q/z2S6yEyHO30XhLIQ2ucrkl7rKNE6+fzSZ9vksGSnYLU7tQ1wUQ8jv
OdFSsqwMwUKlaNSOoUvjaIuIxQ0+nrsy2YdyVq1vKRmampqts4GxbAvmbIFhMSXZ
cPT2hw9ZFJ/ISHRRqgID2IZ3H6QtpjchwJyUemqSn6o4TUR3gscrEM6DxORnQGxi
UINne/L9Z4IwLRbUmJMJ60/z9+LakP8yw4TQSLvB3RNjMuFKcAzXLQxR9FLsz48z
cgMVoc5EN5TAVWdMcguTXNNcJ1d62bVyy3ynEVgBKm58CakqDbxRmdIhTI5uG+bA
Iw5eaFRStRlfnEiqAberyjvoQM6QEW5wafPcu5bKDQandl4B7/xG+LXj9zrEGsWC
jqeugZVoO9CIAEx9xYkGexCHtY4J1ScHzGJsdW0Vi9RrobdkQ4V9hy57W/eU5SRE
4cwgoEzIY4gb1sdIGXf2vJNy8c1RnIeaVBHaNdckul+P/SEpbPmlz/z22LXitfT5
p0FNDMWwpa4K4U7bUCqLMKwQ9Dmhdq1HU7nluTvyjd0gdlHRNtexZfBMOM/dKanT
ybAkgT9EmfITxu6eaHvdyoZdW1KVi5JdB8vWmEzrr/oQ86cMSbhQkUnDQnuhHM7I
ZaUfX11krpsnbkMoWvCpFzQN5P0DP5YmZeofJT0lFtBim7lEerqtIWJdRdQrXjR7
jvpRXEpcLxyvnVnON8yKb1xIuVgJfh6EW51v+xX92MrLVSSwdGiuVdGRh6zLl0fq
bPJYFTdefReH7zr7j1hxKYO7z/qtCoYg2ZYoNyvDLZHP/99jy9smvlivYH3aSbgx
jit27YDvTL01XImB/ItYD5F6oKN/YA5VVHSRTkd0TztOOZoD8HRjoq4xoVgFxB4b
9KeZlASrjuILpeD28fUlMCYZ22PrIxXp+NgUtDlfg5wlu0Ey/DYxdSakDMRb7UCW
/QkHjMFAt0pky8kINpZ9Zy9AERNeK11e0IEyr83T2jky1QN0L85a7x3PKPep7+dn
ag3y5QmTaTzOduwX5c2CTMGfaRvIwXvpTKmZGvV2UDEvnOFgFfjc5QHYGDPWzacm
4uJ7wNnndUrHmYeFAQAUMdtUHhSMs+pWao7/lwhQCK7GRqIzSKxQL4PGpc2I0/Zh
1ECxUHmnVfrhi/CbLRTgfhEOJpxY1XrLPA6V5gUFMdcWZI+cuBUCpPWGvFTbBh7t
M7RVwdF4qs4kytqghmJHmbYwPqg358VqCWLzQU4yfCl7knihIhL1W72fHefRfSSv
mce7j/OCXpg8kRAVPhDZTkLavtzFx3PhTlCxtj1Ssy1ipdI9749h4Jc+Q40TmnAW
tsNWUSCyXteI9Se/hGZY8fU8Eh3xWcTXeURdh0ZXDsvVtaKl/76RNsaVkB2wfWGx
uw2MMQ8NUavecWQIsoAcqSiTws4lDMP4euS6Ne/Fnviduiu0WfYsfHSvt0zdtpRb
BKACy/jt42IaWWLzIZr4Dw/KGnCn618Ah+/iNSr6y0ptIDcv3CH2dG9E7SywMm+o
QcJDzjR4z6EZQed/G2PGwJE0WXHFGM7UGGzKuGo90Z9UJ6JtOzFckjx410SthWS3
yT5s9Tn9aj5q7BLDA2VHEV1OLRk9cGpovkTizD7/WihiAPPPLlbsNezOuo+0Stta
Cb84Eyk1q3Fm8ZoCL4tnB6Vcfm1w4QOoYEFvr3/15sYoc35swvLgXBKigmThrLwE
z+8ov+TUiYjYbtc4x3OIACgmzTkq/TrZvdphIZFUpYwZGKaJBKIvjFjgygTHaS1W
znREdTRbGFKOlX7Qlk2Ijr/pwx+gUxUvYpcaiWTh3sSPmYBteZ0xTs3U996zpkHa
jvmMu3wKI+GiF2Vo0d/alDwNYUBWQeDdS6j+iivo82CiqgiMeK44uvwf4IY5UXWw
nZkTOt9fetBXHfeHm0XLeRNvzoDNwfgnIojPdElgOSFLefN92aENF+27jOzTv7L5
whdW7I5kMAJqCbO4+JtpUiI7dhXVAleZlW9HyNSVxBAyDDuNGn7WxQEndrvuegw7
c+AsxWYkT71yJ3Sr2cY+rxoToWVBRuSe03Ufy4xwzvQUzGYtmz1b3CKBC+wQF3pI
NxVZPsf7+VDUFtDtMzKmyQxqKyfjfM6UzgtaBk4lNv1PFZRShKl6a13YRGUS5LZ/
A5JXp/tNsI4UwBn/cDl2fRpMAbUmyxyeuFTnJ1KqotuvEQZBVmQNqDxzUHhhw+T+
mCaS5AhiNS4L1VW4suXUE0dTMaPoLthK8pTXIjn3AzExYarmbuqXvYmQ4yKcamr4
HEccGQlvW1DQ7zgqKdNUkI7xBZLRIdNOjcZHenBtPTWr/1qIVAlVhlhBG7kvAwJa
yeQv0DggXP5Ik04U1uCaq/xjSSV4PBgxBh4aSP/EvQPO21MixYNJJXOjMlq50a9P
ShF8VeDOcEp2/S0uwKPoWCyly7VqstsSAP/m9ZqcTllCEI6XkrpZfWzr8KnEMv8e
311sgpg5m7C45Kde3oBx9Ec/Kxj2Jiy/+mVh8HJo7oIzHq1mjReHE19SPrKmlGPY
aXW2U0NtYYfQnQRY9PpTi7PMnmwmp+J1iWkXDwEXeitCG4Odi6GfCsz9s47/ddVl
B5w/Mp3S1qWNl1FriPkjrEdSUiGA6lVtHHe9kibOdPqa1P0Pzc6gwiq5O73IHGoG
UACSkPimC3R4B8N2lVIAN8eAlGMLinb4voVron0jnJrPtsjseqd/jp6lpAaOpaCM
vGHT4eq4Ev48ODYq6qG/cPDHuwh0QKbAyLeTKhYlCG/rxqcZyeeS1udvMfeMkpIL
iBA4DRsMl+xmhhOSnwRzxzxOKBwwyJN/euRwkP2Ts/9caqJhlJC6Vxh2/HU3QR6W
ufWS0ibTU4GFsERSqrqw7DcFzJedNI8mpstQqmExtIahxwvKl7vEA7z0wSo46hkK
s9qsTwUEfC7wl6JIFl7Um4Bcvxo8AVrnZEmRv3DI7b1MbbjRiotriRonSiadhY8l
rCAMtIgioRuk+XmjacXWM1tfjd7vyu99rIU2tCEuUAZTjVZAQSmvXc9oXR9lTXTl
dkxjsNvgyfEPtAoWC/UqPNcz2tTdVum2s+Xn6HIznB8vxnnKl3AXWRc6SEX438Tx
xmq5f8eOZULC8L+AVIJldByX6apsegvfsNrkkxPrk0NGiVlpnpb17HGZIKGUbxpG
aC4M5Do+tEQIdxkTEju0lbaciJthBY6JE8M2Af9jK0AsPDH1vLb9ZjrSMy7ijmuL
OpdVtzwU1Bb/nbJO50PMOCILETzT43AkPQ/7GC6H4MktWtulrkJdrRhbF4p7e9D9
0wjrelYpuzxa6DbEJRxHMs0xIkyJLdwl3zpVDIbHonix8hcJwbtbRMfXVx5/HKwX
KFqSyMWYCA0dYbVsQUPC7Dv8qr7jDn9ZDkCbc2fYZ5W/TH8jwAJKcGwoZSAcnHjW
M+iEU8FXu/sITB42eFI32bG6mX6G/R3TxoH8ImnrJno3n13gG16i2zP3NeJm0u6U
+9s/MIVYmyCJiCHk3nGLyepoe50i9deXyRNqQ+RyvTRP/EUocnRi3rOQ0tY89YZg
u4WZnQXRLo/PLUrToKjOfoW0OtrKnsMm0neWhcgEUPjvc44DmlFEBhVFG4RKK/1h
flORt0GN9G2dkf2DvKb1WyRmo1wjPVUZDXrzktlRAn7op979KSA8ve201DSGY96m
Lglhv4rHn/+IL7eb63CHEDnS5V+ZBCQJQWE2Rjf1P83jzyY/AdlnGD+NhDxu4LVG
3kqRGYs4tidlNcrU7ggmcKW3h3vifpUN1gUsF5l04JI115fqySMkILR6pIVJ+GgW
jhfzZPlkT73ypkO5LzMi7NsQZOgTN+6MnauGPbMi/1k/aUt0c8IdfbmtB0n6JMDz
n7JoRQXbiTXbt9Fc1wYhHead2IsDIdMBtYubOksgIQLKjz+E2OTlXpo9QKtjUk3P
Gm1O+H2vKXCR2qBMImn4Dw3qrdM4SQfH1tn7Z0kvdFFFjR9HxvwHi3s6JEPxnTd9
aXZxPO/rWvIMkL5zJRcxeJbJ6qtk4F2X3ZqEwVpNM+hV9s7LQXB+d9/uDYyu9ouw
TdZwq4B6pzXosvUeBX3P5ADLPHjmEKuqU+ZqAavcxdYECj7WuFQVXG3KCqiYrShU
bE09gBv/2JSijg1cm6qyKTgUpQCY/4+jIgBRkBq3kN45D56K7j0Vk+Nel3dtb2e4
CAgFLh79luPsHc5kbcbqcWbAPJQdvEDXDTObtYex1o3J4ltMZX3USCREnf5R/XUp
CcfZpaOEaIK2YiI2ZO58K6D8+lGiozSf3mCzC5eAaHxHjiObNtsNQwGWZb2ZFIVu
tMt8Qj8WFBNfeKiSxOKDYWXLDGjulsXBzR7ZC3hI7rOJAPrUUXoUEIDxeVGAJp/Y
lk/u40Q+zAmz/JxYTt3CZe4PNPtEbOVn1O0h1hAuvyTeqnDqpjhTWpfvmgAtutIz
232e7exs1E/DgtDJ/PVcbkpI6CNFcZR3nljzyWeiNiAZgkimucyHwNiR+FVG4oKS
5WqfCQBKZqxLzW22Zc6pqgdXMlSO5WXT6duGI83Y5tc/ZzzKqGSDmfx/M/CRutC6
4n/AOUeb6mVrunIfIAJnrEtn31WxyZymCkZASHi28uGuOwLJodSfjFMLk5ZDFXzP
ffxMzIQ4jU4BvWKP0ONg0+0vnfoeJvsHY0K/4P6WK6R8zd906lszakFRnjT5RTmX
T0dSWhucZBGGofDml6byf3hBtG/pP5lDfFwZKfIMibaaAf3ZOE6K6PaywfPpe6Dm
6rNM8sxUlSOlSNlF6Ljg7XdHj7ovgt+vqFzmOzrPTSpFV8ty5/2Vz6azEWA41iUJ
m0YNUPxYT3dwu8Zzg6WXTaqNGgh8fk/iMSp3nD3KJ/2D/hSYYOzT+xaHX27bl/Js
izC7QmfPryWHZ8DmgcqIBa//VXlGSmMBvv234Tg8rl9PIqVVYJ75NITOvavWsJFQ
KjyBkuyNAT5iyTAPoQTZtwbi3NSzglapmiTM8N9ig53xUUukgrvoCkY5mRsCkcmY
AABSj+iUEGJIy5YZ2dr1dSzvxbaNxCkgcEfPkbL/FoeiNXNrJ8pZeSsfAkPQgQeX
Bvcx1GcUsxpW9y/Ucep2cEZbN6vd6M/OvNTGiwI4LbhYPvWEl7xWgjzjNVK67z7/
o2Pk9iNzaKOrwBDw+Hrc5dUe8+Ixw2tKm7lk/UEjrfpo5ZB70Y8hu5THepfX3qS0
5tb8il0GLPPBojvDYqxSZYNecJKaLNp0VGc+0UA2aSA9TySdjXQUvv7wnna3XCQY
EWdZecW0Yk8+UJ5ho04sUokxjUymayJMqK4e0wH3660L0JMbhAL1IhAfnU7m8crV
f3xctc/aJaMtxrVc1nPf8wByoE/SAEo7D1K309h5JohHoSS8MzrPtS4Lhb+6HrlF
JpopoivWM+n68KpWES84mHfBDxjJHpqsO/O5rDNS3ve7zvfqynsl7dnR2HrMFl5y
LhAGIZJKXJ/Ld0cvrBYvxzlEvtySyK1XI1XCrvZkI7fYZXlSv2re08dgQCmTkQ6r
7kakoW1MwA4oOQmcAZxCmSthapPRUaUG+3CT72o4QDnXy4b+xbwk4djJT44OP7dN
jSZj2UJcHqNV2CWr0XkT5ZcGZpZilD41H7cgqEKFg4Q/597fFpHSBR4LxZyojANs
CAvFK0eJvOy/6ZzhRoydtNhdCiu/VNBgRTXZmHY1M2XNSKMQJ7DAERYCMmkUqgCy
HAhiZ5EtlNsxWs67foKkPp/JkblwxQp4zRRLnLIa0z7pMcwxdhKe2lb3lcrXBEaZ
+eKIpbSn4ZxoMiEYas2tPsfl489nzSVGZnXXT+uy9wgqMXdF4Y+9TDA3eP4CUqnb
BCZpUULf9P614nOxx7vKY5faBVNu1FEuZxbU0eZwH6cPVU7D/NuE4M+raNpQXWc8
1+XXnIhWdz9kP8kN4G0M1Bl42KOnlHvLfhJrsWFcNA9x26Cgzh8t0+gZSxNmYHxQ
zwvQ9bjAUz0sBBqARKGuDheea0mueIy01y4Km3U92FCMfDmi3pNeLxLJvoHURFDK
X5yLH04Is5g9Zc2GIgEooMVUa1Q8fzGqer9N6PDPLTXl/qCk//sZl+bxIBzRFxT8
i9MY1qCIaP0SLckyCroFafdw8XYHUnZV4Wb8HGnX5nG/b9sl4VbNsGmV4qkaQ3t5
HYt28OQrQokV/CH4rhjZhyerenXQwKaCBO1cZT+5t6M+/CVc123ZSmTMsmveM/ph
+rVp7ScxpkKr3Aw3SXjOdf3GKgDosYn/4AEyrClySJxjjJYP9uIzf9P4LiQlI1hK
QUHac3UB8Efgdk276XvovyQyYJKhASw+2StifqCjSA6gn7wzuXFs5wmVjwVl9cWl
VAGTvemS77dnKcp8I1W3MNfayRUdl4SvVFGgFbNDahGVletWSyqD/X5fajZPecsM
/+a2zB5o5/J4nfIOqibTw86Y0k0zbg/OqmJox5QuV1w9ePXVE51w81Zzb88xSYTz
iPrCi67jC0rie6fCouOVAmQgWvA8LdI5Zrrdx7pTOmKFrsKNFx7++3AiD6jzpN09
KVU0luZvO/8mfibtEzaYYWXGYEmb++//eLeQed5x8ljig0u6g2Ve5WjBcBK2w9my
n381rfDb3TyL7vR98Ufj5kiad4ec7dU78pIYqIlJnAw6bnMZx5GHtyyhZIDz5pei
PCRyIsmJJq8DTFDlLk+HoGDVJPpiz7rILvqxROAmS6RJOZaCQ4ckmp4Ivd9Ksp/Q
mJM1AgX4DKvcVH1RvbYG6BVDj5JU8i+GpKYmiSVpLAGEZNzk4dJVQRBbiRGmywHi
9AdMt51ZBR9RfV7de869hTMXyyD62CWpcbPv4LR6S7/pe6YCLYC8NpaQbL58A6kD
NYhy8XJOL4/BUMMNHENs71wUyyegxfMWZvkHFnGytuYWvf5qLrm1KWH8xkA1HD0p
u/w9fikYykLhk3VrjRSML/tLiKlpa+7GOu4z76fWycLbFJbcs28SYtptBErTv0QQ
YYLWZqBRFBU4XRP+WdhJppFXvzGUutGu3uxba3GUHk9LtfnlO0LxExgbrfYtx89Q
laFg+aVH41FYe/eIZCvhgdyIm+UskU3LWgvqpiEoI+RMRWqNhGnE2tbWudV75ISA
LC+xSTXbuujutS3beRdDSLug7xY6mCyrZYPQzB/QxbNDZYQkEkzefHLy9/1KAOfT
VtstOLJ3GC5QGSWNLLR55IZwn7iNsNjkH3Q9j1R7qC05F9d4bLAf1t8aDGl1hlXt
M/SS3gj8eH8T1Yorri0tj6xO4haoCKMoi/Nuh6cF9RmBSWGuJg35hE2b7IItiFH9
2x+iSvQ+6q27WZJXIhQT/AY6vb1Ei95zN1775PwvZBiaD+OeYG/hA9cJylkl2LWr
a/9VxyOXxldLtraEFN/1YkDWXEsV8krGT7AyS0a69fOgKW5SCLIlQtlByebLNVkK
sEtb2971PTMrwrX03szVgnyUD0fcfKpQpk2FGdMNbt+5gd66hyoHTRDBMjoIn6t3
JOB0PvJAmOcA2Pkw49ZBP8zFHp46HHV72JiX24zQpXU6osP4oOX383vCChbZ7IBp
Q0giZFIHgjG7GwXKFT5TBgqQst2I6IMFR2LHKBzqRrwViHN0SPpabnXTB4ib24K4
FSjr+7Gulb5CImjlpfC/Nqu3M+F7gkXkLVmo5NMubl51ODdvAVPtTwal/U1rNCIB
HAwgqPwua72yAXJzO5eAqa7Zxl2UsLnev2qgtg88sZw7t+1o/bwVaOZo8pFnlMG/
Y7lE89xAyqSRwStbnOciIh9JG8YcQOdcRtGzLWK4dZ7wilyGn0F2dOL4RiCJ3FcW
PNJrFFiQ4wkvYSIlqBaFndk6P/+kqXpFTo5yeLFmiwta1NOzOaV4J1QoPQOVO90H
JRp+ys/vjYK4DdKsAXGg1QMZ/qvnDwf1HMctx8u3Csv/z2/U6OKZT9ldAGt37aIx
kkOnzTtcE1MTjjmE6TTwNXVCzgHLlpbAxltqySVfeHXJa+G3O/DQDlBEXG27VPJA
Bq5hWAiQwZ4YKHt45oH7a4RlTQ4K1vB+IiUJAgSL3M+jNMbcaY7U1YGiXni9os2z
61qLD0MnXvha2fFiaJ2UV2hu8nvtwdW6eZdYQF4P+ku5MmDa7//BjWDXkyufQUul
/DHAW4NAS7nu0BRqj2DSRWRhoWsgBVBUBD+5L/G3YFZvHP2BfIDe1pqk2Ut0pE7x
ShFGDgdI7w0fBKFumSSZUGs7h1Z2pzPMadZyT0M0XY6VCnrWJoVxo5TtV34Mmv4A
U2R54c/Ifprpn0CRHPAkkTdbqMA1yHiCiI52QGVcg19Bt6CzT71mc+JeV7b3IDye
GZr4x4d3J09pjCoOUx+51gjVWmzDiX0EfNKX++p68XfmYjg2jQVP/pJDcimIgLHc
FVe0uA1PGeOb10LJyUBr8XLIwmZAggzvLxsrJBbvXTpMVIX4c2KBf3rlhXgDjkzz
SQJm1q2j0LUCU3CI3gf3nkYtYA/wEi93shJKsEzr9lPVm4BR+KY4Vc+3TmfL2XRB
6KuLaBr6Y4yWNFA3ZXmfBHHr6Yc2wUbx12nG3L3yt1qbtyONwke/hbP0WTzeYoRD
qIlxi77bj+ZQIvbeqjxr5NHm3/cJKVEbX0Z0wuN5zK00SqVmUGjdBiT6pPB+dWba
hG1SPy8cS5hlvgtnm/Dj66iCnW58cinJbvuc/i4fnqQNQLPFIkLexYKWV+bAK9eN
WlDoZY0+8hFNgQRrCcdvygYsfHgTY5rk2a2momk1M199ZiJ/3NAAP/dcBaSI1vau
q1ylDMmyGZdPz0J/fdLCRjqpeDEoE/qgkt0LdihCs/BZugtLIJb0J+dp1pqHW3v3
J/PJJqGZfv+gE3vM4kpiDW2qBJdC9Hj06+oGr5mFlK67KLxGtfV/1jZsM+P0Imm7
a/TVLvjT4VlegsXSCvbCSLmLhAfY7TC8OjYgQwrHVJGPMqPDj4XGFp0QQBEA7+GW
I3fbt19k+AcvydAmiv3xw0m6zIWC8pcQQAxiritdurAfrUBD2LA1+ANSqsNWnj0a
X4MVrha9xC7MQv91b9jod0mPsxBzdhOD+dNQZgIGrpZmW+gfTlXqrmf3rrPIQhOw
/WQRlWzySM9FGJlOK7um2HoB5oCkvA8mJ4VLylcRBr3P0nnJHSkh+wzOU0JZ1MwR
8xPis3yg4Kijfsf0fj1asyAGY/WmiMdI5ABF8EU2IF1rfNRtUpk7HyET7iVuBA90
Gur1VyMmpQ3hl+5qPRMHcYlmmSwABsV29HN7ePe8vrEWx00zGBssxG8DPiLJSofF
tt4kFy6zN3UvTNUNzPmWgjytY634hW6GcpUuK+1wwYyNRIUT3Am7opLlrfP3HoAZ
ZzS95fnjX0sCalBBUv7jDB7wkO2YutSDKx3dH4+GvBKYFaqJWRFh/HD82WqQSvHJ
Mte9aeLl0HtMbVO3pHCOCsMnLeGFdptzlEiJQGSjd+cy3DOe4iqNhlg27OgjlIhZ
dKvv+FZKpfmfi9ObcvpO96NxQ1/tF69qk2EI2VG3bU0Uks7Nvc20qyrfFqXcp7H9
XrOz6qIwfWWj/oiKPbCmDcVNwccqbMVUoxVbsBsI/mC6/0eyjzOqg3C1wNcg7wVP
rjCx80VIpzs14PS3ZSflhgr5WJ27FOkWN+dmx8h0K0Kdd5eM8IL+K8vzsOOE1s3Y
HZ6htxJ9bCB+fQ6q+Exay8Aja8YVRuOlbYcA9MOGBiXeInjVInio7+I9xyLSi6FE
xRJc15u0pMfQsFTGgsAA/g70Er4XwwfGj+F0h0rMLm13UoBJKwsE/riJpdMse1Vd
Cfe+BO+rKLcIDoBmYwgs2vu5ZjGKnCPs8+Pl6wMckhidYGfLhRCYqLgrIbY16EQq
blATRbuWewBucTWm5wGtlj7yU/+FctX2IHLohCFN5aoXlFStTYlTZ28/f+lo3hoA
vtu1+tn7eayzukFCNG+R88DbDbOzTiWVnIilvIZstP+up6kPGqrZ59LH2Lu6X5AT
hCiE+WlwXBJBlk6gNY4/hxavoeveHzyBZDffCF3XxfN1XbS5z03oRmmPiRAocuJF
CDtu2+v4l0jfMwaNsxH1IWRmjFRLVakR77pBDL5Hz4mGz0SuoUEEl6HFUPUtqLnk
oll86VBACwu8BQjZC+1H7Gy1x9d8W0wQs5oFDXmILUWHjK7+zwPBc8NLbJVpYo+a
LD0QAIqdeZ84GcD9zHqLgKmE+x19RkijdmyzqOAV5eSNWbzp3YmhjAjXW+6nAK8U
MTdjqwyQtYXAyv4pqbmOD+jH17Jb29lVTWUmSslCidwbRBRxdlsLILkHmk0lXLbL
vAoMe9xxr60PSfTATC8uG2IsFjklpHBDnlJ4x90ipjDOG0uxLc+E6XmqLIoVfiEY
E79oJu2/LGIu8/6w59BRI5iTyhDnKqWFHculW+ulr9xEp7KMj5qEUkj6OyQmVCAR
eC0nb6PVWebbNwxmNh4+u82OiZIClkadsoXsDcGvpyXXjb7ylfghMR8rrQ8RVJCG
TpCyaIMuf84JV/RQworhDD8kunp2eKe7FOidg48JMHQbZo4lH+CO05OT7WSamAKY
zlBEhBOt5bWEXtWf+rP8RjvbJjH4EAUdIj3iQjdFBE2IgkAyeQlan6Bb8VpBJgbP
tla8dBzd8NemlCPon1wqfXOMxTv77pMY1+L0MpD7Jun08RODzH5FyZT20Xkscm3l
bLLlFAwsmKpyTAdbEu9daO+bI12SvrxzS8jevI6WwFSiVJO9rYMMW/D4E8sunNmv
6G5rick5I2haddyecEgzY6kx9XOYWfskamXYCN9bPBY83PVM5eWRDyEoPkVwwyg9
TGuWeD9LiQG6hisMUu/xP3Du+sxvZ7D43DuWoGv16SgUJyoGTVRAFEYJ2FnVPVlG
Q5eIYncpeOCq0ThounruyCE4QEdEF58QjNBo2+vWphCcc1smZoCcYX/n+2P1EC4j
c/aocDuViqTDXpE+n8rkTgB/GZkox/TOxl9eoB7OpbZVVHdZychznDxWpLDr3Nqv
vJwhQNqj8J9T3+YnkY++XdupSzxeFVOd/Hb9C9s5bPT+/f5bvwf/tFC8oedvmX9H
9XqRMoGUEbYqWAgOJUx9/e3SbnIh2m+ln2IAGTTvnEo9OKwjRihT65uII9e/CDP2
q9wn6E1NszsHjbLwirlcSkqVRGrli+vvEl86cadSfzykQvz463dichM7yaAqCtye
sTnl4ATibltbn8gxlFMsBYHU+K1/8Dm/CiQOqGm/pXqqOfH6geqCFf6ttS8Fvq+I
fYcHFw2aRCayrFtefDdC/x3v/bY99CUILr/0Zbnei7DXvyGT2mzoYfZtd1Ss9vhO
HeOP9lrRmrWSxD0acJJfeDIRrOxAflrsRAchXpXtGdk3ri9PFETJqFwSS/Zro+p5
JgPviGgg+aj99iwqr3fRYth86BBK/OzqbJCPMj90wyhVXc7Cxi5SvYHXRn1zF2ZS
Qwz48OdKyoyRSQlRmNW7c4rZ1LLYyvnRkJ+vDalPVHl5wITJUrITqEhDMLNf0IPc
xoGGRYBvS0GOLbYF86BdDeqFenPc1mqrv/t/MSldnKHgPmJQCiyAoNx52hgkXLeC
m+tiBQto4KyJP52uGigIfCVezt0ZWAC86eNOPB0XUW40aGaoVy7YyaG8R2bTlUPa
xQQJiITUOKRf144taQI/rIQp2XyLn3PRReHt06a0fIT0Xb/eZMPq+zig2j0Jr+zb
0Mj3f+yuMSU2MqvnboN5mWAQ7tGjNP+5oBfpltM9tWbdTHOYeQMYCJdb7OfkUHBO
9u3AvD9qpfkMda18/jWdyx3yHzRnA7c/t0HUhmhwr7l2bHoZNBZOSdOsfvjKXUwj
ZbnNt+Ay18ZvEeAR/j30mFYlYwbKMx6eN1qF0UmAP8epDHVGJhbx2JUhuPOaovbo
mtAk0z04gWppLbrglrsNtCoEjjfphinVwUJn83tV5jl3MssimSgoPh4/tMS3oD66
97MsKd7Bz2l7FlUDqewrhkLIXXcz3Gh3sm/DmrSeuFu9OUzr4J/RBbv048U3yeVQ
0vw9qreBGORaWz6N6J2Ck9NVzP5TeLmuNv8pVOMZjF0+cH0r0tAD0BPGZFnwuWV+
5HNNQ4fbEGNd8dqy4NBzJ8aFaZ5+zTC0GX4O31kEPgAZAc/VNs+QN6Ij5LnSV+cX
aSo8qtt3Crwd791I2QLeVMiK5BFRqtXr83fhgZUvLrH43mx+LJH9DfxFalMPX6fx
o/tE0qQ1VDw1vGk8/BN6zIlg3RpeeawrraAfmQXv1xqlpsB/z3CAYCGa9TNa27YE
QN+7YKG4XZ8hHz8VsfDRk2dSwL+hRnLiYnvMJPf7XLTqKAOgxhjC8IQFCcGalW6L
PnOvahLY1/l03oyBK7jA1ySek6qbPTGOC4JtgOmw08hAsAj3lgfgMxL/V1yFjkxy
qQbDDkzFs0Awgos+vCdtrnJOruOjvSjXW28RuYuiBkheT5P2BkX1mcvX8ka26WyO
NhgZdcA4wF5HmPWzLeC87v6yEwT6Tg3QzYwgEEsiNGXu53vp3HEq0+ausNVHfBs7
k+gHi+86J/wK36TnBYqVNKQXtTx/D/rIh9b07fnFS7V7TXCHVzMq8NwRkgijRYwX
xHR8nKy6wHAVI1WdQAJ2kgqTDmkDHfCqUvF/3iWRmVPIuGSVajX3QqzpMrmuLDmQ
eYPSBFU38hYvVZTcKYmFI+jBApPJGkfH21u+i5IAEngW2JbBCwqg/tJ3m1+sS0VD
FgcdPfH2hfGLDQaQ111MsYVbCUcOLOsUtGiUDmcLyjYLn/UwEzf8N4vJCk7mcbRq
Jt7k4Uribt+MIQL3P9ZAPw7TTe/hhzkEEAFFsnQNbP0W5po7P80bvtzrrY/xz+Tj
dNuFOKCbmPkE9cbNRbW4TeyS/ix1STCZjDtmeMnt7+NOjV3quLgGMC4WkdWiIyuG
kD7oQRSkcQ1K9J/UEp7vdITVqiATyZve8BQhESBxF9ejGJgD5cHZ7BbGEtp2H3Rf
yWysGlRThJvhoxhi4C6Q/8MpcdaA3xdvyv90VZvraf6VZvgDtpgTyJGqj00JHFGt
TEeImk+2n7XLrjJQOjanWvUJuGdTe0kFpXw7Gtv8bhdEho1//2wPYCjv1NnE8OY5
b0OTHbSk7v21r/Ppp2e5EIXLWf5kNORa+D1tTAKBouZAUZCAJKaLVLe88YUmDmck
PGRiY25oLJijvQ23aCoRrAZb9QJRnu2J/WgZpojBT+lXKfqg09fNEyKdXCUC5Ebh
RPr96UHIVBjG2c8GUGG+1OsIEgUgRUflu63sfMIxCkjuiWhvydPwgSEyiC0vVUTP
B07jNEIwimRwGzgk2mNjSyftLQHn8xgi2xsKM1oAjEQqCzt8gzCfmW5QocGIQOkF
kP/DGkgtbsRspso35Xm0sYgrdNaw4XMmi4Oh7K+s2TUHzpOTHHEKCau3KO9oZ8fl
2+rhVoTU6yFeX6va0KeK0+G8wDA5gAkmRWhONzDbu351/an/yQa4+oYIU91bhhwd
HHEAFsTkec0G2B7o4Ipe7IfTRgORLOLz6jr3fsnhf+MDRVvvOUW8aSXKLrEl6IW3
N1dbDehQ1CP/tvr4//8OmMqMvlbmcDPoxSDbbSR9s8nWduhp0+7ibI+Lg7sayRt8
49TiBTj9SeNTCbZ8mSVdisHtBk0KINmgpI5tJE66XXgIaGNvIxmB0Ipumv0ML9gC
uncYpoM/Wy7k9yxwuf9rUuSycQoYBSeMT7Sef0pDEzOq3nx7Kb2ifeh6Rtva3XzA
sDHjnhpl7YiT83BOGv9CH1hjzFAl8BwmcoLGBVNOtTKpLMNhz4gifLRK9PmmosH0
vuWtnJF5ZE0RxTaNYqX+Lh52TDce8Aj9GIp2/pBXWOwXTtInenYgriT4f02He2wD
rqeFX2DA/GXc3aPN0jo0xdOOApL2ACRhYF3WIJRRfIXBHEhekOmnL55PnllNiOvk
f0l+yZXhad/hdvOMuPLQpHJ/uTywoK1H4r9iZhed0S3t3YCVjLgciVSkQb/1F8qM
qax2FeeVecPdLd/kB3BWEtei/EUwFf2UVkha2XD0f9jsBtpyGb/gLAFPzqvNl3Ld
P9RNYq7cNyawWGj5hnOIodUP+WtselJA2cXkLE9h7aOZE5jXxXwEZLRwLaFCaNpR
O5+E9NTx8B7TaXxWHkAWOC0qk/zRM1kk9dpoyEWaKfLGR8IiyG6lS6r2X5sUrqaA
RoH8Y/g7s87GDecdYwkTJunnRMpyoo4pjgiH5BQPEfT0XzSC+c4gyUqoseSh8FLh
TZq7EFGTAPuSFV4NYPJOyconyzzruqQd+KC3QXM0Xu1mfGFPzxK4oiVMY2oY2ACY
l4Fl86sQkITZMPhCdHit22k8YdlnFyeGrdKjZuSnG/pzHQYpatTECDHADzG1mA+/
eLwpe7YzTjciqMAFYgE6EpLbzm7q6pca8BQygZvBC2Hj33O9IY9QPZyRfUoN7WGv
/1sBS2vDQe0lsdYbcuUKlD8fcwToxjWyAneJs9IZndIF37/HRx76kDma9BW2vXXZ
vZQbvV5X14bFwA/HyUbddyX1DA4VC+AXaHzB8WNxMdt5QShLnKkqbtlxdPtX0Jgb
31/TrtY0nftX0OS7f0dtQafKDp5Qvlt8AD3NTsvvQra/AKs2vO3EzM+60orxIA6w
6KbrDFpgL1uenjUHDj5L0Yk+G9FdwjNBkPM05cU6acuwCZk5HH4HXLFpiyurhBWg
p6PabIKmVv1RzM8eXYK4IRFtbIQBp3vVOr/pUtHy4SK4+pbn5qc6oBLt5PiKy7kk
5u2W+MUrFOpki77T58n1zQOJgoeFDaeIsdeaAWGSUeI7LYjEkQtxfGvaH+Pack7G
k9IV8038la8wc3yb15wyu+3BpGUSxjDXaO4S6wWps7ayNf+XfuNloF6bXmpxO1qi
qJ3Lap2SY1/45jKF0oLfa59GxkMcujAILfAxAbADSpsc+X5XTG9PqkJOjFJUKNaS
dJsTPASsGRdgXchIRb1OjSR91uiga1bNJ4u4siTYim4QZlanM7Q0rzIiyAW1Euw6
Et1Ha3Idmu2g9JoMZ3RlH1K9VGW5lSKyT6PKEdy1MkI3gh6aiABCH+RBNk5A1dHk
vA56rcV+ANGd5hyeOEg7GqKOjDPADYmLlldTAQa7e0dJrvoPDRVwAntA2WGBqqlm
tg1j6ERfxx0t0ne7KqS5Dg==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
jhhm38qlX1lXoDCT3MtnBCZa4QKUQeOZnn6qbH7f0HOngztCGrxucsIlt1cDOYi1
PlH+kw5k4e+R2miqjFDFdGfvdePAip6n7T2VwyITaDtgdxyPnu4ukTSTofh1eZUO
eATbXF6E3n6W0f2gHfA94TExbt2W/X9n1voXpvg9tUs8rzxlxYYpfOOBZbSVKTJ4
PMHy5aDfEj9+9qx9hqMEnLv/KxHYnArn8CotUHeB9um65bbn5TBdHrI7kFMcGVQ0
VMtvj3K7gQkQIomDxuwApu1TZ9BhN+oXbocNVMA96IVnuHYNV6qD50+8yiiVme7S
rByB6WTz/HnyylkyV+cMhQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2384 )
`pragma protect data_block
v7CH3o287R9XXDjh8FiYL2VUEW5j/qmUKRozxUhr//O+sbSiUALedfOM7ZnF4YcK
v8Yh9w4tXxGFIXUgN9iHV3JGJiwzyKfbUk9l4MADccze0HKHVYb3BPFgp02Hqvvy
2dHxzHJEDy7QopfVjHN8bLvDksJgaYV6KkhzEixx6XgLV2V0he5uYgk/T+Af/5uS
LDS28HiL6vZLVLsdxfX1WFWElom2rUFc74fDa4uSg2ifVd7Fm6Us5hckeS3OydVd
ZJHgmaBZIs0fhunkKVtOcF5jFcSWNCJRlntAKFHgRzsFyol2j6tH7X+tIoAQPjIE
g7ZnpSwD3pvuRDqaf8PsiSDjKNkPtX9QaXyGh6HKUpFmDTRKEMgL5ytqyLiayciI
PAx3oCjflcVfIVlt3W4MVKfnQBjeaSr/iQ1dJpyCBBbqFYxGz2lww9zs02q9fvK4
ItPpMc4qakxny9RXuIGXVds8ZhbJkrb8TsAmSyppqae1+DFIYcZUinQYYOOSPZzv
lOnoSuOXK52R/DlPynpg8tib5P26ihbUTmykz77JuXSxM1FdUVnsIcLwMqvmJeJC
Cwbg54Ezhu2wiowMO8US5AypVnrBT0rpULdeAg49ejM+Cx9+wKLBe5Ip8hoaGIe5
iD3JAnKi+YYUSpPYZHD/64r0J8QQVPOgknVvsSs8pUdukZAPuPvkC3I8bQg12apq
y9//G3GEdNjUgRK9RlaHIwEPFlON/ts1i6MHjLkbsXfsHnIuhbnDqZCDwrWSHORY
2/CQ+eX8cL1gBavES6YLePqMUC9/GV+v4bsTRfQdbcI0qxViUbOfsoM+/is8uhxZ
p/OGeBtMvtRf7fdAQhJfPZDRFuFHI3ccQpooQJfGTHPOLL0CuLcs+QjLrDNfKibJ
dZeX3mDmEykxyGYm+H3q2IamiQ7mjrcSDuyhk0ogimapFwXTkLvGuKGviQtgjvAx
zHLZvC3O9xpZtnUZVhdCjgHUU0ypAfPiGjl4QfrdHcL0M/0BiSM6kpXYxhNK7XUE
e/rD7vp0RXxUoaw+DDo9KKH4rFCfsbUjcMN2B1KBGx7O0nr9Ip646kuleaZqG835
XnqkfBIDfN06ftcjgs4vQiSVHtZqikpB7eYSdQ8yOIKwKIuxZSmITily3gszmM6n
eDol1TXgnDbA58jY5YPvI3AuFMYqm10ZpaQWuRykcOf1Y+dH2Mv7t91yQa5T1wLJ
pN1mK/ZHsVKahmkMnLbZV1jrPyjiOyBaR4vDCYAWhk+rs161eoptlx1dnhN8uwNX
tf5S4Gqj/Y10Wx7CuTUMznCXvmpOK6Z2AuAujT/E5+d46oqOd+jjankt7qsd3//B
Wl2WXBLRSWDlcy0Sv07iK+5889ZpOPb6CH6XGfbZzlL4Ctd2TYysJja/La1jQPL5
AlEU71Boio5p2KxSTMgOR+NmNOVY4QPvwCUNH1vINvj2RWp/48hzoZm9XRTHsKFU
aOOhlb8AMEU5Gw6H1Lq8w+mSKwyqIHsS3IEXz2JQzVvMjqhVKp4vHBb5SqPDx0oK
Rr2Z5IXWb5dKUpK4PuUOxOB56vwquUJKYtQrOGedI2Sijq5SH8/yo7Zdxktnl5JU
sj0okbjwQdAE/hIriVzRcCpt+HO20QUJLhlKMLS9EpeIkFu8WgeHnfyPomE3MzCJ
kEceDzuPIcoOaJpR1reypiHz861W/q9MoBetsLC1FzcQ9XFeglK4seQhCWFXZG4b
aHc6Nacckzjnlg59FJ3WtfQMz+kiyc0qfmczZGk0oCOGDMYCWcqQSqpXsdPnts53
nVCt5LInfHwPjo1ZyzN9+HPsDxPXed/qRI9g88yyupof8U0+IjRtDJb5Rot5yVAt
d+F4QJmKMIBTqs2Rp3opJzsxjp2mqV7Tlne0+lqGUQ5DRDJT7XwSqdIchMl8qm42
+4q+ufiGQVFHQGaGZpinMy0rkWh111/ww0LpWSVGo8P+q1wBdDLFISvfhW0YEIIe
BH3plVxA7JN+xkqcv56jJgLK1i8A0WqgUA2XtbxMR2Rd26beLuMpMC/ctAYXo6wY
vAAHl2tHAmO7cevJ2VguJ6BrUGR3Zc4Csgue5EBgfrJvcHW1S1HjvU19y/mB+ix8
FNlnwqJ00kvySgdy8A00ROGTXscbGtbh8bAPZATrFF4h0Qe4OBVKiVXpnet1MIpR
WzCQg6d6HaAi+xzw6zw+7g/LGl8ENuMV3nRNaW1I2/KLmUKJEDkxstcy4R4nvS/i
4C5iOSiL/mVyXZrg/eIOouIFJm4QL93hMhdKMwIf5r4RDdnTMlqT5f47XAZ69rIU
5CgZhyuvZOzHt8k8WAHYfrzKM253wXg2WYs0q7ouEFFTwlK7r9M2CDUqCcJRdr7P
IXJPvwCWFp6tZH+8y16YTkS/IctlarBO3vUsQ+s87f7Wx424ug0Wlmf3xjfkNpkj
Dj+HZt07kEtd3ZVSY0V9rnxNG/7DvRbgsPxZlqbOJRc1eA5j1uaCI/uqPQoYx0Pg
kfNHIyzQwcxS7bAoWUw0KNYitVwIxXyFQwSoso4URaK0FKdS/xkQdhyU/Y7SstyK
J5KEVchfakvq0zIr63YwUqdPcH/qKJ/O0rlnIzZOasoV/bMo9Qmz7QN5ahB4QkfX
r9XN27NXb7MAwx0bCkQD6Idcf5DZjiQPaRHr9hjHyo2QMMvrt5J9dTw08kPdLUnA
kwUi/1Qkcuo2b0hRgbK3LLs7WNH0ffo319RpDkleyJuInbygzXnq9D8FLj+fjXYF
e8Z6jhgupOJLyX0ao+8LeC4/xQRsOZ5pvFR941hOtQjPdz/q+JM+TYcH+ODPvU/4
YJb9D/QAWu6ryO/H5+m0f83gcfLb0LLfR+6s9fnuczEjRi3AncOnMCuOjUA/8xZb
bP6HTfbrn5rIJLJ30KQd7H8AhwOHF2qTGnbCs/Faen7Nhx83k818qnsTDuwueb6/
7VOXggi3+AqrWrMvgF5w3rV50jpFpVyt69qRKHfXiFLS0ZA4P3T5m1ZSm/ipvyk/
FwK/W0I2Stm4E3eb138HSLtJI7Y8FyKI6dp9Gk4Nox4jO6huSl14kMp4C3fw/oVO
BXrpR7eWGDUqt09Vy/5jgZuJ3B+uB+VYkwO7Je1p4fUUoDeS3AkeCBz4ZAc01qJG
4DFVpLxvhSxyoJxzfYypiP7vcmwrsmvCSZnpn3BSiAY=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
aVfUY9SXjmBfpFeuBs3COutA8an6Zhyias1TZda2NH9nf4LGUIJ9vBKLFUtd0lki
FejbPMy0R1rGWkkwsg08kdNxjnCl2PEc7N5V/MSITBv99RhL+sNzUv/S1Hlq2xdY
puYBzsZ3reyygre0uQg2aR+Rdu+jwUixuHHNYB+Y7/wHaBsv/hxQzRHjDtt4hiYq
zUaRK/t68CC9xz6JTTjQEXM6ADKHUg/Iv2O/4ElYnQpdSov3+UYbkRdAOaFgqnc+
uCQqxDIWIz8241G6eOa65o/xS21JR9OnQgqpWYkFV7LfBxM//jVkN/L9AOaHzVIP
KqLBTOIMBZRulyoVrb5Ayw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9360 )
`pragma protect data_block
712i8dOcl97D0CSVHB8P2U0XKTxQPZfjLVCKppyRGnWuGl4UXiXEq7g2xpgcLZR+
r5LMupYr1qm6EQqTTmwvqrYcOfApTt99dwO6u9Dy5djHzsiezIZ/L9WDoLKHrIAZ
ty/qCHF4nWcsdks+obLRP1caZtrv8SKhIP+VZBvnG+eov6s6ExeZuArYJoZ5/CFV
PSK2RoolJoNWqAqSfbu+M5NihVlLjQSLiuYIg13DkoRVbWkDGw/mOy5MDyCr62Fq
sAfFy+v3Jkj7RrnOshdOBB4eVEJFRQIo0SmTWa4qdgq1sIBRkgTeycXDVsgHDr+V
JP+ERUx6tNnGW6Haf/BnIiFTWZfhwdxd4ScI7+aGe4xwwUOfzdP8V29MYeLjsTyx
0DEO5KxlabeZVRyFmFV7qpCGg2q9UVhaxfRLZMinop8I3SaqgFwTAFCRxI3K0wJ0
QhY80ccFSYaV+1pHmgBzJBCJIN6Q6lRNe+foqc3zZS9NfHYlTCXcHnH6vUHRNXkA
A0A70Xv/+u/6gklozt0gFQXr7uTX24A2aAnyCZfgicaW1dM4WJA9GCYyTdg301A3
YUMH/O0GeuiyJHkohA1JsfnUvKozREYt02RjjqsFVoFLa9wN0I3XjjBrJ6QuS/pT
9q5ECx26P/O8WVeIqFjT03ruP5B9mdwo02NCBDvn6AWw7Mz4h3pFODFpmswthq9s
XIZ2FZEwdja9ZF0dSt7f9usVCsAG5uI38NPe8dsCLskOoL1z47JKAWYay5Dw07YO
xr6xlX3cQD7En1h/7zgdWgGoEPbPB4Vek1fm48NorkrndroxqKtBBd596YAgFgHh
MNl1RRxvMmK/iL80QwzFlq29xtEDgcsfiBcZhk4EINenMj9IIVoziPdGx/anfCqA
MOaRCXWup33e2k2es5/Oq4EEGNVA/q4/emmU60o5utAGTTP8UaiwkM6zbCvNkftI
Tpgj0+H4o97qPJICR0xjU2I/oj4PVlRLo/eR02gLdZOo4NFPEHPbYvyLJEPAJg0z
ISka4EDfktMaufcpZ4Q4JuUPtqo0r7ubXvPVIJzFqNjWXhOIGG5anTRU1kynuLcC
A93KH8FT2xI5WBFgn/dkbqNmS4db3UbaZNuFYKdrKG+wdX5qItrcEPJ45fKLLAxb
YVse/WWZAt1BhMvGaQPXD2dyOOQvLkl7amQ6NEEv/KLF3Fs/up00eiF6LSVf1Jk3
Ck1xSFcJz66cOrNbecNGx9Kbgx8PTQ6vbUtFT9bijIjOswp++nFnpod+pBm4eMOz
PAtJwRE/piASZ/1yvOP23bd5raNvqAUD17v/rwurbszTlfsgZ4agWSk7QY/SBV/F
fE00bONrs482QShWnOh0e2R9c+AxFyOHnwIEiPXnasIQTP2knTRTFLuyA7cJoemf
Dr9P7X+XDzzPsimPVylktjBrV3HcZH+yaqQWfQLTu9dbiXpwKYMKr+ZK2j96yNcE
V7tCTZUfy81ZunfzqR9UWbxpKs+ZPbHy1P76UgIFLgiBLSqYYrNqyGesa7NCfoUL
o3VW9i9t7WBnMkaJSfYzLAu6Og+63R1NZFTbSS+UgMLjbl5yfgqEFSH0mdu6MGTl
GbYVYH1HP7I6cw5Q4kbwkoU5cgjtG6y1Hqh0SXqCZaRZGJKeEtrofZOtZXTvedJE
O5ENrrRLCqPP6nfOIgXKb2l8crs1nhF4vhMozlDiE25sLrG0wF4qA4dqn4FyMhha
mqPveHZ3vtk0DXppM4at+e4vn0JEs36x0Ax9up0uLsuEKZA4+4hozAPdGnKG9KIH
SUQAKqk5G4eQkt0gRnlNFCmv1W8iFIPnNWK+lu+zfYaU0hkMkMd9nOc7p4gHDQy9
SLzI4XDEEEl23xjYvMM7x05Ysj2EC0cjzqjCk7VIeFo3/cP8NCNkZCdsEobeEiyr
OTtTkesOcOb76Ead5nUpaVyIMClqQJ+sD0RagnTC5Zug4v97+RevfwVIJE9wZhuy
SZb3b9U2x46To0wWg8fF4Q/u6RIkJ5/rvKrR0zmuve5nBveE8gTssrx5wk46j8y6
PEWpvOEtT0wxMIT9jfqVNpO/jZGMzrj7k+0EsECCkPwjvMRHTA6QfhLcpsdx94D7
AzKkscLtlWC6NWjlOylnPCoQnI/7GC7dULfeHlgqFwSpHGLJX4kQtN+S1ifBcapn
YHMp4qKwfU1mRXgxweNGanUu8Am+tCIylJBMpVpir2JKw7PEDzSvBe39QYjcTznD
+ctt+UAwQaF9f+lbbv7izkpDaDowXAMiRxR/JOFwMIzMz5fbodMHndk3fDsifH00
PcsCUzYQ1V9Z6qA0NcAywxlnwE69OvndFMwu0nMSs94D84hDjUJ58bK9gQkidgzX
zXwGMd4qwsULSi9BSXa9OnhNkc67poNH+8tW0yvJfRuwE0bpRPZ2K1ALqwB+ljxA
YP5BGNC/5wAODugvteIzUoNqBnSVoB/rGn3S9Ro+WyEiX3kUAFbD7cvrdhJsjwRL
PavDAQjNmtaHY6iBkOdSsQnwwXjGUA2fni/tqZ/K0EEXU6ubCPEM/9zeOvW0y6dg
NsEFWADv+LRDx9V+nmxpTM/26Puj2rKufTMSsAyIT9ad1vfhRvP89SU/IYacq0f4
D4B2TL6KYKDw54urbr3zC+h0vcUlryrlfPeq+Uiy9kuO9BlXEDNE/TUEJ5ceuuP9
QXvMlwtvgKxYwKFBq1srdkKOCbO2bN19cWbIr59Es+zN1llGKEfWN0dkl1mFP9l+
gWHPoW0bI1oRM7KCGydOT+fl0srkqD80dK9/r+GeNcEKj6N9tzvQVlVAhEQ1ha9v
Ypn76jGqNkbTGIjK/lz3EoxH48Su6YSUNXLYnRKxwGPhcrVBt/VAQfKSGedlYX3o
Xlm5qHfw0f72C0Qvlj/mUxq87PI5i/HfR7N1yjwyWedoKkykH+dTgrULile0O15X
oYmg3L0I4V0Gc39o8crWm2QSZsaV/c45vRAYi+c7RqFdksdwEmkWtkRGs5mHA0NC
yekRKS0DQ+Dz5lZNw+10o8Mds/bv3RKpstHHBqHAkMIUs6hcf/rrTt4RgSAuqvzs
S1M4sUMY9LFMbMSsYSWIFmPC/NK/+GIvruTeBQPAgO9bE5VV8y5RDO17r+qlPzU+
1HikgDye38UJizoXsEUhgDhDMZrcBmIBm/31SK4m6ofhNLjdsZyTfgbDd3ZCz3p/
XRRMa94j319jtcFJwiPwQKyuHFQ09ubTday1vbaDK610whTiYSdWv3DYqsKN6kc2
LMTH78IDlVWqdaWg+utCJtwu5IOszJUOZNFK59xBD0gZvCgx2Oizyupe9DW9eAtD
meyMF/rUTTFqAsmx6SQCac9TpPy/mI05xdOj7syXcE2j1GkCdL2Z8tgT5TlNSdqk
XeuTs4a+0KF8mxaXTMTbump2BuwY6BW9fO22Jz9HlpW3UsE4lfKIYzoSPPZMYqMt
9qpofCa40yIIVLljYxguWIDSoc42TFO/xv+DoF5W8xrh1U2GZ8BkJfORYXXMBkeI
OL9sVRPPgsBR5omuyiQq1MBUkasnzmg6Bmdw7Dj+K6geR2koyqH15dJxcB5F+e/P
UxUE6tjsOPWikXIqeiXW+9ZJ1gfFtMK7R+9r1IO+Nb8I7MzVilVG0oLmk1I79Lyd
TcOqJQBIKBTAnb4VBoA2nI55d174769UkWK/iGs7udFvznCf5koAN56hbt+AC+4F
9WFajCX7VXJJqB1zuC7pHzoEO2Hl9sRj40L1Ma6CtJUFXzfGlhIyo4PY1F4NK7T9
8CGRZ954xY69BdueWxtr8+ukUPK8lUx7RWAvg8vNmOHWXbG5xyzoV1Y1DnagMmWU
SGF/eXHmaCn+eITNiVOXacQi3qJ6GMXwbZyZBFx7p9sy27hoqZF7tlDxPLoD9lb5
QOdzLnF2hZDV1cW8s6JQQZWSFExdPvjhefS/aga9d9hYkRPNcbFM0HMk9iAkI624
gaLMtu8oFaGnzvoiPXmzQKNkB42OKW1sT8okLC9Jlgiv1HGHepr5CaZ6p+3jB+A6
FS37fwKyf2U2xVbVFrVgvvPFBAdhA+g5OBYs6jFFZqhfbkNOFbCVr4Swmxi4Ntzu
cwB1PS5T6ZYzcnZ7p3z/xaVH/QNyXv/e8CnuuWN9yskFClV+axDAZQtikkWHoh/4
T7EuJjJg+NjWkG9d8DfBwa6gZ2/BRwHXbAEszbh2rj5c/Rmgz5KGx+U8I2qQ9Vgl
gdOsakrwd9fWbZ6UXGIom7mfD+gQqe0ZWdAeAWmt877ALmC5YsrnKPhiRYS9yyN+
NnjAhKgXQ7k9NU/5gmBaRyI5J64rYmyDMFRpuxhgC6DzfZaixAxfS3fje6A9+nGJ
I2R++QWA4vzFJtw79oFE0TWePVriWS0oizAjLOfIZJyWEOU4V2AlBEbhkwOmYgJi
U3yY546v51gUeHGQYWDt5SLJTlNuI/XUEXCuir0l0Rhxu1273UmJusJ2M6HBGqxf
EsSsMrwe7kXTvGwMUxRI2WLgHkYzdKlnMZGtJZUyuNszg1Vm/bnk6IQNq/uArVnB
zbuEvKRuJ//z5Nw8AfePAbHy+krV8aoI8SZgxykgXASwY6juayaHvOdKsQwCDCzX
9pmhF65LDJ5VdWZ2nKYzMDX6lShUHDanAsyhsaH3o6mYV9xi9aSEzD+JOXLkp8Po
R9+Iwjgb8FJ3f1vEDTS9P3u1mt6teLkQZV/JcgEkZgLZZCNd6PiTTD/Rbi/V/uMl
Grk0tlUBMApseKLHYvhJVWExuhH47GImYXlH0Xjtw/f9Beuz9SHw3gQp6+dJvqm6
seeYgAetrCnxAmRVhaQw2lmTsttOOPFeggotHdPJSQ4O+vS1BQDqx28ccT1O0QIq
GDYj3CTuGEPAH0Ke5RupnhyGAiSxJgZLLJNAZFXWGz8rDlCFybey4FPwt6QS7Ljd
TrVJK6m6XmsZD5t9UnE0XJ0vGSrThQL5Gktdpvq2O5gJA6jz32uHoDm8AEwt54lK
D9pvBLmJYdTxA8FxD9NeQmpkYYzfhhEOWLmV4tzY/VvFwzofgLENtgBOgzl1Q8XH
cDy86V9QYMtJz+Egd54wuJcgmz6CPQy/XC3AL6h4z8QTzqZ9b1yzBDXTJI+SqbUP
Th0WTln7KI0Alr4p7ytAPAsK+B2/G5zQXqaspVKj/OkS90HmcZtTFFw2Ya6LVVFX
4QSCdonPufWs5/kdPiYUeuZ1PefCS78z2HCzPzJL09HTmgHPzIS7QrbRJA2Q4Zdn
l5giOXgqiBHZm3GHetd6Q9gMt/pHpxr75Ux6GZWaRziS3Dnw908Bqq4sYvW9sqwo
qSJGyoPAOxLpTqQKWS0i5t31TDbdbvozpWwev4f5e2Z4+N3PFfVJzQmli5PHjuFl
05+4D3NR0c5QoPxEF1dfk7po3NJITOoA6jGVPv4jyxWyz8FsNuZyaKgUqJXQw8hz
uILIHt+vaYaTpps2QMSJQX6MT81wD6YHCUGe/IkAwl9lrodYm9wh6F1Ni1wsMdB7
HcfOYbp7WPlVdLmZy4jcYbpIbVcbpwJzH+f3PsdnH6nlSxuXiYIiMG737TqPeFq8
5t2c7njMD0Lf5iWzqfZrqE5okMH4a0zjEKRO/o8mURxdGhzmJqWuZ/+/O5cov+nN
5HclANNXgiK9BIX0r/8dMBycQxLiliAKKm5TVkvug1q8W8xDE6If8xmlgWTYJuUf
iNvu3Byt489peLPaqv8yPa4wv0rIfvIpii/0o4g83Bw5L8NIQLqCtj2xqpwba3wX
RAGkoC0SVptfrUBWMRNNK6QCklPuGLFVsFlssFrY5zjv14LJz5Zgt97UynQy5wZT
8slRCRGyYvMnQMJKmrIyppjR0VKjPcbYYupzkQeNqfewOD5l0SzrLBntIo/HbUmS
Af6B+RqpqmS7OyFCZz1siDrq0baJPNTcIA3Hg6LdE9jbkze/S4oJyjUlgBEc4pY/
o0DffJaU14cjDz6jLDEy/OJm9pSRaJuRX6nr8UxFPKsPvBnZ9jhi9sJy+w8lA6Wi
6klpt+x2PKsLSk4hsFMJCX/I0tQzb7RwrEtZTX75cnVwH9ANgctBpdH6LSKPjLvx
+9RRmBWOB1Z3Vt+5ynUFDyo0WzJWAILye8XSPu5PjLzKap8uVGwsI0i2uKOb+Bg6
Asp+YO/4JPkj5fqIGMPzede3Ft441IqVHDHfFKOfRh3gA5FRK9F9TsWh1Zo181or
iC2jyqymNTphfyZMkpf0s0ZToQZCSQd1fkGk2Cd5LYv1LNLHutLboq71csBEDdEX
XvGwz+0h66s9VdrjUSv4ypWtijEnc11+aWmQKmCRaPIO6DL0C092JOTGC1XQ14QU
UDs3WRVJsFBwMvIVSK35RSpgEXRqwfAAiLvZYod+seSeUrVBx2bt5s0IH84lCo3S
prGE9f9EpmyAG5ehk1Esx0EVoBkrDeufXUAVoFc3siX8KvxfnIDSg4QLGPOf/j0N
/xu1KsP0gThffhJtx4uVjkneOBPvfnLNXDqEC4NHli71NQM5VkV+LJLVO435iDTx
ELMnImMVCNWX7ljSg01CKGQVkLnjeGlGg81hplr7P3JqgE72ZjMscwnrsdAvRNCX
htioDi045bI6E7a4Wd4Pm3NYWRSJ3GWFdtnF4qsd/b3FE41jqosaLIUFlK4BG4fo
wKHHKWt+TtjBP/Oe70PwumikOqIOOIif8JJ/hAWfNA/B485uzOiP+YJH9lScE7da
WXY+GuauWA5xWVfMsqyV4ClFiJKsfa6Jv4L3n0tnu+6IZWmsAotsuQDAXT/0cp3x
B6xP//vCPZ7vbbKbIcosX4aJxD+nEkM2XnAO+NqbTKfMsuubJNXaA4+R5qyETG5p
hzhB2LgCpI2BGcupz8wqHPITaJM5s7uNUOCMkGJyRCz9YbSesqZNNyYa1kJw7S9F
D43Kw+CJVg2mHTgLZBgvePIZjCMoKv17PhD7Jsagv+pOKSs02/RauKN0ELd2EMIN
R5BnCDILfRv6zeFtfSohPwNtBEjJVgLlNc2Hu1hpQ2Co7YY9chWaZbCyp7Zt2XLp
J1Yu14Wk7epUmITDQX7VKM1dhdLgHHJxiDueJFARI2V5zkdgejzNTlgWuAt3yvCd
1vB9rPTRN18WiTeflBZQ8JLdWf9FbYdP3BOHoxjy/sikc5BAuwGXhW6wPQfSroBW
cayiEpKM362N2Wjofv2byhAvXGCp+AEmNwjtPXZ1Hml1FDt0FFP211uuOiyYnJIz
UBbmoESeTk04pBGIeYWHczGkSpC3XScwvbb8YmECgC2j5GG7uekPqZg7Q12ZOulw
K4R41UvPDdiyYT6alF/Dxm5gB681lo0XJ1jN0AxCZjXvCb6BHcrSkHur9CRNPCv9
r5+qAK9Kghg/yxxKBnyt4swKgpRce5y3sYNcLluprdkJDW4B8m9tF39Z+iHAj/xV
/btFjq3DHECEjydteQXaKyDQUd/Tww86kWTQ4v4S+KOL1j0v+38l/Cq3lf9XC0nA
+BxOcv16IIXyJ0pcwBKZOWDttLzLOyEJR6ixtlMXHQbnu0aJFE/ouwejLEgtsUby
eY3fx/OwvET/kRJQQ2OdHQ9AmeIIx2TDtEqQfMzQe1d/GBcOxxFf9EpShtPEgkNG
7yXDJb3Q85B6dTGMiPdhHd+ptZuBDz51BkvUqjueCj0RAwvVZzE1kS7c4CjNApBv
VGr92Bdvz1Y1RK2xTPDYENfXWqJqkL5xCMXCypKo/SoVr7w2C7p/Ga/ehwBgTfq0
/JKThxLAcTvFwF4a9BcQOZAoG+ttuX1PLbweK2Dq5CEro4uhKC7SKt+rrnVdgXx8
Rw1210boFxMSKC3jrRt91AbUZrRicxDGl3krLRqgkUkblUY0ogfKjO6maWayHswE
u6CS8yL60QuGYwL8qWI+HiOYZhnBUE7io3+MBAImd//eK4zsqcqyD7icFtpjJe59
eoJ/M/ath7bXvBOhKwYLC5sgEueHZOHv1vCYvNSY2kmuYzATf9WkCtLJMTDSkVjZ
HtCrwfRhBrMcMqduqqBA7qsOGqOMjfnbF/kWSWPyk3JicOxogWv8TdYGX1fUCf/+
wvFihidFkdwAwTRyiaYfGPhIWgwdhFBlIbhfJECu4QkaX6Gd8lSuK1gs8L86L975
cyf2QM9qUxXisV+fwtsEGiDVuSX1mDDbTuckECa66KDhl697Zx3Xn9rcoOkeV0NS
b8H95i8SbwSNP9zQ6yGbhr0yrurQq0c90KunwXGZS/TG2eQyp4aKD57IRaRB9Mh2
0NdouyQ71hjw/iYfBxrypHuLwUNGrUPZi7AgcmvHfNru+JhCa3Dy/fjm7jk/roSq
x01MS4ttowO8CYA4ZXj8gR2XK/4rm18JazTJWXi7HEn9oP6QnJpG7i+CoxrcSbo0
HTikMqbQhuYiGwLoz9HHbsVwzQzRjb/TctYkAQxiM4XjmKW3deHMXKMdAnzqDgUX
nbfm3rSzLokL0MUvO7zhv1Up9944I/hBdbvXJcRpRfKbQdTxo0FxfvXyb3LeL/eO
r5JxOIrN5rJlI7CMWUYE5t2wJSgMHbNX6ryjKslY6ax+cT8aiw3q+BbfWnmItznf
4uUjs1ukJs34yCEOYIG61eDEZQ2aL4MmRE3zw1DFoDzjRqfzqZdzNzoEb/amrArS
IKDZ0WUKgM13y2GLWa7SAJbvn4PBQ3oB23gAnB0gfa+YZKjqGKLrHy/ANqZxEYj+
2lx5UhL4/NfWaU+MP+9JEyPlJzDR9OLfYxIGPWiYaWjcFd/fCgKCGReuoNIC5IWT
UHQNIsKyYmDY7XwRVpXCDv2617MfIx17CCqtP2ecZSYuJEG400CN6A1bCFm1hnMT
yU4yjf9GjpMMc17zLuv1RCyKww5qsf2KuOtqtFrhRa9bLjQh0O0KHsTMRaeuueZM
1mwvr1Hb/Z8r0NX4FZfpenZcTv2nEUA8NGORfNvY2AuFzYS6fsFPU6Bt4/yt7W4a
5n+bkuuIIEyZ0xMnLVn5HKC+bK5lga1xsJ1wTVp1lRuq19Hul9GHQ3VDsnCTPPVY
RSNKA8i9zRWChZnA717JCHDS1VanRqbkXsftp2SJbH5K82cyZJ7uwX8s8giudRkt
3NyJ9jj+5WcDVh8USSdqDEIxM11FwP1AX2QoVNEC1yE9myIIbLf+m5s1XBD34h1y
SZP8JEhHO4KHuZHTMIbqX7y8p4cGahxMF3jguzf58otO8UtPYbrvLb0OYQOOBy3F
bwgx5Qb9tzOSXQ1ejnFSogMis9QIzx4USH89Dxuz1Mm6bbcazC18yNuk24+aJT+m
XrYkRK6xvWyHsrB4OzT07diHfCObFqkQx3zy4zDPf6BNhjUxReUkOQiNJaVFRPY9
9LXBMoJtpSveg6geEAdYou5e0GODpKP48jnOn5spB6EnAwREtbZgbsM+Y7D3H4B9
fcjbbtxWHKM2TXtoZrzXXy+YPmakfcxyI8t7syDECkoDuBxhQlckiKn1+eEqhMAV
bUstC4cI0GC1KgmGFhMW2RXAdEt/IAOufU6sSXyNI5vc0TbU/s6Xl2GoYlkqczD+
oPSwHSWjySFlakGqoL95DJufLvQsUWESJaPY4JsxXyUz+GzASZpHSgcDJpLsrBJ2
s/U7Zhca6dKwERRsE2EswvW3YWLOomVu0xkssmKDVE2L038XGiK3CsQzZG34HJZS
acjGTz3BY2243t8t2VOi3D8feCSgmuNZJarDQwRUrCHXkJRHFeGN4z4jWAiqHzO3
36iFWu2lW/5SgoqzTYUYnRIAgcH4wzQWH7y/P3zKlKhnrpSvzlA0m4aD2NBi6fns
xte1l/j1ny/XvKIv5CIdAo7isppgxCq9D/9eqiL2dqEsa6s4A14IuisC3rgpNF2G
QQnEbaWNXUiXZGXKQ1zA+w0er/2SfYR/IvL7GehszEOLYWiTXVmwV371pevoPxL9
78f/3n5vAnus3ivP1VRZ5QnNpvKhTJo/kSQu0hs8LnuwfcEh/6iWcYWPxTMab7Vi
/5+j2jeP7RugZUE7j62QI3XnUNn3F+SMsfScd5CDk+08mTugk95mtj4FaB/BFOVI
C+Vvd2H1PnoJfEz9YaQG3cL50Wyt71D+1m8LKTggwXui+dW4RUQW/U4/4UPz7UU1
dwVlTXWO9PMZTvAjexc10cMH4aecnjiaMJXmfK+0LBN/MizZ7yHqAqlNRTZ/msOb
8//VkQKJ6RGX6FIW3WGXGhBMPiDeSjCydtjnnYPpd5w2uk8ybZVDEvo/6xIT49ZG
5rN4TRVZbfwJegGH8Ln85gt13jAO7ucnyM4960ap4vRro5WNJCuWwUA4itVwuOMb
CBWFugSvX07kXhewHocJ4XhTIhsgtUlUitkWLsFEqAeVUTDP/KWfuGCTXkJpaA5P
ZnFh7Sf81cyxwwiz0HWVh8VB86HXxKOs8Sj1UGiunqSoSx2rwe8nJrJcbQvj6cPl
/IHKUHqSTfDaz8VINu/HIBMlZGRRMQw9z0f69FSaP6fCv9NXGmzjLy+uoWJJX33n
KBziaYWdIPq8hJ8m9fr6VgH4DzmL2dqn9Jm0ZQ9qClW41ykg3wjjbRlJFIdZMTaA
xJJJS8KSXGlU/Xmxsff8op51jRdK7S1B8Ga+FkGjSvXCuP09rNsbudlAuNzorHOA
RkFQCNIfBncWwK1XdAFw9a7L7XPh3qjCII9YZGQjWq26Fe2lMv+Mpsxg3MeP6oDf
q/oSyo78INDmp5p1Dp1Rx2OjuUN4y6ergA5w4q9tu25XwUQnCPIo7D0P0AwvaRCR
4d7ov47Bq1kjRLQ6AWEZH7t39eux0+sQ/MMcVTb08WpUDGy/81Q26vwcMmv5tjEH
PirY27IjAFC4Q8QmA6DnI4KREEGg7VC02X0fmEqT99/BQ2zw3czdu/PralJT0iCb
gD4ZQnrMZExh0Q2Bqo1AywUQyOJCApIqtIm2Ocn1mYzBkutLwHugCQaKt2nt1WNX
lZa1EtieT3t3+kR7E8pRY7mrcrV8Qkw4jEuBiYmiEkXYIZ2DnxdVj1ojrB7GqFOv
dNnEr+39FYzvgUYQg7oRadhEcGs757CcoMszKIz3Od+8cgYTbgQjpLL9dw+lI1Fc
WCSeBbch6XJbVQwKUcV3TkGWeAp3zCbhI7wvJZ9QqkKRm2x8i5sV+8U5q+6lCz8y
/zALA+9p9/aGk1r6/SPPBmySwVYhdcHgb1HMKrsk3162u1WPaBBzW5SntnNxm/IL
EsEDauOxcF4utmvpv5tyEFwD9210x5IFSkgul0Rtvw187qMXu2A2wbslrzTVoroj
2gncKeYduRj69BSkn1z+FTAQgaELs+jHw88xXcgo/ET3aFO7+DJUzGi0kIbVCNXD
No08pm7ZHnBmiCMU/NJhMAg+ebBjDz79VIKJq0ff4MoQAWeZnGLLv5dZBGeJYzo2
K2ChShKnpDaO6YW5IffqNkG8nByPw608oTBMK3Ye/ft2Vd3w7tRmuGXKl01xFIH6
9M9tYVY7cWcCnvp6USSQUf0qmZLG9bWniM7e5zrB9RF9wmkUjkQWLoUC0++1aRZS
It2KMyONKmP3Vs7j52qbNfVDusASgonjpueqlHIm5itxPHVC4M2V/d6WDb62oeRQ
h2pAg+LnDoMkr2uaN7la4QQAsHnFvu/L7FEnYfSwgyqEjUejUGMpf3ObE72cr9yP
8tRkfNV+DZBz36gTUpN32UomsyuLKaYq1G5WmNiXib8xVdxqqpiT/WTJ96MERPWu
Iw0tEVetModIavdZWqr8YGzha23XAwHRd+se0WH+5abA64PuomGh2ox9mrG8MMMN
WyVpLplTLzVJJwk1x8/X6v3wyawHcXB62pE6MvuweTvY/XYA/bZELkr7jvzmurXR
irzx+e4UaOWcJRI3VDr/0zduacOQEcHoNpF7gAXv6JJHtka/daakkeV7bfY9epic
aUzrvyoC/Sra9GWnCoCXQmYl36KW9tOCYxhlt00sjNryIdmeOJl7jGtw1pd+iOKe
YCz/73Ik3PImGSoyDCJIr8gaeVDGMR6+6RFPXIGUFeocaQC/HLvhfnAmgMgujLPX
8wlinRqlAkd0P+D7Jch+JEYop36nPqBgcymXv0wAWSGH5jXjXjfZQk1GOqOAniPc
LslcLp6sxSgonQwulgFLn5ou9WDbHbEWioA9LDVmDEGntZXTK9Zz2ZpXj+UInwi0
ks8T4R/AkTWi2dh2weDeR/lgpGTcOq6uaG5BRtP/YP0OyXjf13ixqZudg8/AWsI3
gjHHx5fGOkna3eo+hJiNlHcj+xa9S66EB2h1ENPV3dxVAOl83hkQzhXqdpU6/iZZ
9k4N6Ep4+mI+polX57RBzEq0wgR2K5j9/NhzrAxj2FEa+A/VgS9yJLuRAB7I+atN
LMnmIUzRjy9A32fD/id6oIOfW927Gt+WJRl51jAuVJXdMtko33C7OxP7BGFMtnmi
hfZAWTkGp96rTGOgGFBd6Om9kk6eRvswaDohibrDDG3fGXFqiLtg5ms7kd4TMho4
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JJcfu0ktzr8u6UjidmPzik2mHDOMpIzS37I+JfRsq7BvnTFpoX04GJYdsc9hQVYk
hr6iTYi18z1vlx7YzXAPV2tZUvS4HYap5QqjkJW/S+fOAeyOwFcXPRIlyo5EOuYM
28j2Tiyd6GIuWx067wznmjhRMO/y2fHtyVa4OuoVpXM2Dzw96WC/wg3mngfAI1Ns
HK4YTrhaptUYwtawtKoPzkyjLNX50Ld9oZ0D54VV2jcZy9dpM2yYDP4xxb3oXcsM
X34PJBPvbkBbHxn2koX1r94lXhVIfu14jykwtjM3yJhG3QOyEOWczRyinlCSydzS
vb5+7sxusqkfnwoLfTUhbw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4800 )
`pragma protect data_block
7/uaO5DtVD35BC7lnPdlhWq5U5bR73vj9+uc9ndJFcBRttI+bHnu+2WHwhAG+Bnz
DHMVdrY0BcJXXJmRrfTGcFJQ3YC2p4sQtmb93MDe/D/6xxpSbxRKnCjTWV+TLRO2
hEnICoXbJ8Pefpnmwcr23GPLoRmTrsOa6cxQFlvSivyOddGQJNiFjwgTIlgB0x4h
Qp4qZ3nxz5ny8RjIZoe6Zl44/GiYBfylx+xZtVD2mG2MuqK/H1dhzE2RgGSyrQ+Y
CP8zGVhtujM7KvxZyQZvNkFiq2lRONyV5wRKUo4Ff3YlTHnEv48kfJaDUic7klRA
Z1w7Z2LzCIrZUcfbO49/Pj9tHkP8k2LeYDOlqsWKvGYwflz7YydvzY6EvSJSK5WE
ondienF2oODWqz8q/IIEsBpCckeG102o9IMuZVlhxIPb2JoJZXK7gU5kTmYG9gnT
uY0cIdu2GxST6bgdyYcJ4Uz0VU3EADAHPJjt4qNabvfMsfie6J9aGJ+osceiobyT
ZyjojdWSKGEFiWg0TkqgbDtMYwj19+A9QvmhddNuiKqMieRQWzueelIFdIofGxQ8
qxZ8yGstpVyU14uyd0Vwl9LjT8hGlyt4E1X6+x+PMzEljMj+Nyxp34QNIo10NGOj
jHuTDjcOOAr7g2IphdtsKQQQ7Wcn+tyq5LMU3T8R3q2hpw2r8cHGPzSgp0Ujl/rs
+iIXzaVt+td88+budj+Vs52TTMvauHkiructAcx010XSh04S5+dgPQo8bBJeIDnv
2TqU5NOD6YTTc1TWJSyKhJLLIQIwzZScD15Uj3wlH2jHJ4o2edV50wme73uvKJdh
Ags+Hf6QF4m2Z+KVa/8fzbk5uj8Gy/C8hhGdDosntLTanJ4oBGivUQyQHNg1Iudp
kt2AI73wBrJa50SfhqqHFICgfzQqBD/BRnaCeYtqLioN1Jd4VFzhgCncUwLReARB
3ANKszPe+D1JjLtLV5sPwoMFTcCJyHQ6UMgBjCtQ+uS2dngKFWADw5qNWGnuoUP0
gXIPBE5EIUVbnoUvAQvaMFA8y8t1oAlfGV6dzcWJSb225kBiOT9IqdrOCpZBL+8v
Yn2EqUGekkax9Zzi4l3IcVtGoDn9wuL9W4Zkq4+irytZYJRpFI6cHS0NivY81aS3
xtn4/fRlFkjmT7zkHLPAoJbNai7sUpI7Yg7avjUmNXuiv1m8lkTk607b6S7DvalX
ZfoHsBhu6IULf1R8yZ4lYfjCSSaZdusBs9FGfGDLjy53rgqs+T95u/if+d1206gZ
sbWdAmqgrX/o2qwoE35gm9ietJdeYMjNOH5IvA2Vj72NJSnBraacxFkLIQOAPyll
TXRj2OxD5BS6SgD7kPu/k8rspVrrXYkNKI0PEubQ7RtAyW5sVPpZX/PyLHIKs4OV
eKLJq+WyEOPof4g1Kt6dX+XvYgZZ6pi0bBmZk9QdZJWCKaUDa2Zh2dkBnc0K8xi0
q8IDtZspN3qixQyFyQqlZtSHVNvtV/JFcoz/+4jCxrtH6zXA6bNPh5DwWgm8RxZG
P9543Av1JZaca+MJPTAghUyb2iK5uRp7Q3Jl/ObMzDNaLRNtVGWnLd3VESbwt7Ut
mW9wHISsvBq5TMkP1/p3vyKUwcy+QlFEqDSLM+goBbQnZjHD2nH0VBaXXKIo+UfP
DvPCEwnPsYmGkyUyzIRqEb2rXGDKQfS5+9AaJvfKiWp35iEsf5YIHLokJ0xUsI0G
lqr7GeDfkmnlbA15wW7XHkypJkDZ8At2EdaAGBJELaBbbH9gywnyO05mjO/NQJuL
zKFpZiuO9wn88y5v552yv/XXUXylvq7PZ4OUn4y07VbpOlayLHM6nuv1gkHgaGhl
XvG82IoqSAfzrzXCFY2dupa3mHXtAAinIkM58ko7N4hKzkmuEUXg2g5bvcY84Y+E
vVyIdkCu+8jwg4lxmQLNTcJ/vVTr5MfsuxpsClvy6NOenzvovnJig7itacHk5hEQ
LSn0TQhOTUkTpL5v+RGe4TR6xZsAYTAcztvMRGvN0pddrwkOzDcbCIiOoHNCxD8P
/BzAMGS+RKOlj96ItMuxjOMSPFuqWaJTPXrO/u0U2GvTHnoz+1q2Zgdm6vACtAzD
U/oeLrOeL3t/1ACKisuT8ruIXLagpT6dI+d2satQeFoXBocRqsjqHjIzB1U5m6A8
1fQWGU/WZL1mtHEjPatWiMra/sQh7iXnqJeQWonlD1uKlH3W52djSkJLhBSAZ5B9
VoU9YT5Vc8oaFlTrDh91XSC9lh3KCwYO9bU1dCJdNNEIa/EnCgM4/VUe2+B+GHcv
Zjak21UK70KEZvGllN+1ezbkxDFmTcn31jRzSWLvbN68FuRFS3qUIdF3a1nCHgr2
jPHf9BFkeHFiuOItXACQKziskk44JFmV0CVLMEGTgX+jRofi2u1f4X26MGVosmzR
ooJXRQTcgZady/+NQSDVtRa/R23or6pfRVf/byA7mKvSs+SaeB/FFwevg8ul0Ves
ABOTxYeRE21Bx/NlhroMvwTNLQHwgLR57r3axCG+CtQYNI5QQIkfVlRVyo34JZGc
39rDW82s6n119ntIgwuWxp5FxavcAsK6s/HrGxK24CY0evyvS7OhnD4fDWBwI4/1
Ziw2o2v3YxfZ0CXGBscZ2rPEOt0dDO/xNEg+BulsBFGs+S3DOItQj1l/xd4NUF+t
IbeF4QOsZhZrKMAm5MsOC7Db+1cqpf3VlksvymtS7aprK14U6ECnstO8uQiSPNpq
WVtNq8mRpYni42DJmMptSrrQvDLQhADKW6jU3/Zlj8zXxQPpCa63IggA6j29g0QG
sW2Sx7qjcgc8rEGiXJxGusreSWg0gAdtKPkxhArU6wigt8J55Fvt7kAwmTGtzJCE
HfpR600sWp5WVRwEwp5/wpM+hclMa63PmdaZ+uNzlt8QE7f3bUhSD37CyKvzZT0H
o/m7KK0vHqdUN5nTqtge3bP9nCMa4qnVzkJ2D9VHOsC+FFrCqIJMQDcj6YKijZ2Q
YZsFa0tLXkn13yzEAq/r8APAZ1Ca6Z62JKKdy8OA/PD9v3bVA6AATgKLO55SPSgx
IIyw29QJnridRTBefe2asCjcu+SqLNLXif1DoM1Vv67T/WBIosvccqAeeP0YJ1+3
cwNjoyi6CJscwuqci4MFiE4bmsiVwMDp2dSEumZqMlNR+9QBJDR9GfdgL+plNu3z
wYciGTp7yeh94xKMnDYQr4RNnCTA0RyJ6VxQKLZw0e+KBpnBdPsNSBtQF6lPc/AX
rpToubRfioUGiwrJrGznWq0qGM6vcB1N3V0WUnGqMpM3kqdFkAQQc3zWeA6HLuzk
pw2Hf/oaCfYOWJnd5LSPmTdqjI7I9fn2GdyV0+2zzu/1KKGQ5eGkkNPSM15d92Me
Nq/GgnjskIOSqSXOr4VbygX5J3/KvxYF0W+Z6Wt+o5Y1CmafyEXg53qWjRwE6HWW
9jpkqdaGmOt1Qinoux1gLZMrjv0O+SpfRP5VYPH/aa/RXWmPbzEIafsWasDk2h25
oI28EBXeS9G0vwcl8dBAE2kY1HgSQNu2Kj5evokkYk/ZaqCAEl63XnuVhF8KdHvA
74p3/EbhQA4nh/llk7gGRJ/w9VBHg2ocyeNCvvAitomw3iYnblMlbk+D0m3CFq8H
S7UzW2yk3Aq3eXFm6Y6FrnUI5IAebIyDFM36FZaL9KRu18BP9QYTzxB2tUQtZIWO
DaW6mZ7FbvA3vqy5KqyDScaYzhlzerCL/Y6o7FkSznAEzjf5kDpatq6yi4E4bET5
TCeOvwgYCXT4CfaxWh+651CxF66TBJV6wRlt7ExDk+Wk6GNLO/BYBp71YioCKJl+
UHlct7SBBSc0/LgrZ3iMNQMZMY4xHVIE6nhWIv1Wm1fwD18qvHhHUoTBZklpI5Bo
KQy1H6wGS+0zP3uDBnD+iPLGDiIb1mIowl4cA3t97gB0wlS8liGEeiNaDPazXu26
CV0Tro/BwQNbV6CtVF0UOlxY7m7NBfOoyrykPGl1bw+k3bN1kfIE8Fub1RkEQe7j
n+dr982bAd/97VqiTYdsP/Pwy8mQuA6dsXPiko5VtgOFhJK9pG0pnLMfxdGHx/ni
OMPyMnNo1hi5h7nZNcPRQoYIAg9+GSFPJU5mZPTkh9WeUfdrPAa7ifaOoEcdNZFf
gfht3BMggxkKhv7GJVW4WvxJr1PeRdsA81QOL0ITd43PoG6Fv3ed+7mAvmXkc4oH
LvmYo8km4k1JtFDpTpH4J4u833e1g8WtF3lKgwghhpJsF4K9nFB0zp6AfzIrvacX
RB0szj8pHtcL5PC/pHymov6s76LBc9c+riVv/0vMEKyaQo8eWPIvnDmwuvF2QRgP
xjtV6ENE11LTeib/9zcsXwVrb9LSZICNzP7tTXQ+2EYlZ8BMAhmiPpmw4qVZc9a1
RG/FHQy/T8eiS4XlzAD4RfAB1FLJG+/gzCdPp1ZXRELXCX7vEG6GhTFGpRZGGJxL
t8r6NslI8O1vKqaqu6GVoLBFPPbxqyO4n/+IyhaSK1ML9RzgTabe14Ertvj3rP7H
tXrS43joaQFQYHWAAVMVTaNwu9+22RV2ShMOBmLhL+SGx70/8v58lrGtBrDIBCA7
BTDggPTi+dyIKscx5mfkP26kYamvnKqJKLI9SKqz2Bto9nR3tOWxlYBoGbGQ2WUC
DYkQTv1v+zqOdmjoJeW48OpVOja5N3dLZP+1LG06HPAf2yaiCiuP5TH/QpHJU0VU
oNJYpAMQkKFwgZhzdjhGmxy9Bgoyt4/YkQZi28rAsahZNlZ0lCQXb6tt2g28v4BM
Z60wQPhrOGL2ePubobUucvKmELe90G3sHV+0q3C+dy/PxXZNzpQWmMqHpjxju9fw
usqt4H9GcGTh1mQGdjBvXE7PH8xdLVUD3lxN/BjmAU/FwvXtzCrERQgePcVWe/wz
PQ6Uwqd6NdpuBRNsu+ZKSQ58soG+Oy4F9F7Rm3CcnLmkxKYkV1ym3bBfiiiYpD/G
9/uLhIia83VHnnKrwl9S9KtpYkx62kQebAOrGHvgEVe76wQEQAAcrbG0Sh9yHgu5
uoRZ+aURgCmAXcL9/UliGC48JQfMuswBRo9W+sjTRJW3Lgyz5L9Cu7mHVLTLuhd4
4+UElhyltyrjV0kXjz6aMn25hjhLz6Af0L79FvsJasCxTxHgD+6ooWN2OEbSz3HJ
tvDulnVqRdjfJMEuFnGRYaplaWiziXhTXNj9zmM4xP24pKNEldd1l980BL7qFv2V
TvtdHubRHatA4XVttrK/I5v/3usdUeEfQqExYvUFvZMAdLZilfAQKd1PN7r9iNWz
KtWBSKUwLPHnzCfO530vmZ1YQl0fq9z6xEHpeaTgQ1zy7ElSCY0wB48W5WISwl8j
CQ+0tRMD6wMAvoWeHOm92Nv7xXJsjbCgKNgoY4H12zefZhE8Bm44YXpw2dgvOaq1
E4VW0Ed8oTiPGIgu+S2Zv9ShsmVTyHXkRJ6PlvWaco8AG56XtzGPhAn8/yBc03wr
uNXX60un29tivoLeDnF8cduvucqYp9SkraNztmCQPHX6zFXHNmNcSRLZcbwJyOCd
wZu7zrxiRgcgUzbkjVaKJp4j13ffQY5sQIONGJ4bpakE5qbrkHZ7oNjOKrHu33LZ
3BaVzxGMm4qNN2a8vw1v6UHc611pKFgw7Af/x0SqMYkHjlqi79nfkv236flT9SVw
rDrGjcu36L5OpkKXQxZkB5jnBp4vJc2I1wXG4slIbLuQ+Y+o/xRH7yDPkLHyev6H
Xtrn5gegL5+u9jGrM7n6GoH1FVbyGZJWaYc7V2PIoHouXCyCkSE8UYnEgQsvwQRn
p18PntUFMJYNENRL/q37W+0D9xyQmX2R6ACdoFGssBO6V4fEFUUgSdkRyyzQkE3k
qLYH9kaeZdOFjAUZjgj0cN6mVE2WHySk7drd5VrZCoF6YiY3n1uO9GVyTQnMgBPh
wj3Cux8kP8Mrm5M60xhfSza9v1sW6Kfp+n/oMWYVoSl++EGQucyRXYdlXNKE9dH9
M4Q0Fxqv4CwRlDYcaMxJwBt5dF7xMzho5VWEsaaiM+PAbJhi530/2e+Tvx6JplFI
30XS8q4OolkkPO3RcKNz/0PqWBatT9+Z0hjovqQ3cG9oHqccTCF3Ln523AAtWL42
NpRPNuU1lcSJsAvAf6HMNn3cwEuc7ipNcTwaWUtngD2U/c4GsK/i27hpVczhWKbp
sYOdxuxZFpvg9TcDDvtaYzJanv+Jo3z2LqhQxdu+FWmJEpQNhxflOQZlj5Hkjfw6
fNtG2UlwaycLz1d118u0FMnz6Ddb5ArkTdcnrQMYM4fm8T0CtpwYWuQIL8vTQAtM
/xpTp4AUOTWkkdxVteE81SvZsgdaLOwfIHolB6qYq4m0dsG/BKQXXF65rldQXq8e
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
KYxJmwZY1djNdPXgUM6v7tlENk5L012lC54n6LCts7NCjaSmhM82XQv3pfjyaw/b
47qmT7fISOHfhlDXkj4wpjRu3kdLLanj8YEKcwytb1v839ibIsMIqit9trffqgbD
XzKK86L3VubmXpZCBB7KrggUiJ6riH720W9AcorTMNh5PDJPma+2GP/rVTHC/6hA
cJLuWOIyDzXJlwlAQ1tuo0rVN0ntzgd2OuI4ueaF3NrnV0t1dSedaVJ50ksk0x9l
PsV1mn+gC1B9sd2gcdPSbtR3WJ9lbpY/gJby0+RY8AcLApIO6zE788mMyU2n1nSQ
3Qv2MHjo8L3ko3b+ruODCQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7344 )
`pragma protect data_block
R/JDIBjyQwrv5WIts5xOYcpujw6RYgo00l/EnjZQIpFm8DiG+WYC5W765tWYFWt/
pYBjg0RwW7UK98x2E9dWdh0JOhAknQbYxx5svbnkGKgY0lkZjssYJm3pkAjOq1e2
+AuZ2vcNS8IsxS6efCm4V/EYTvoNjjTX/jVLwUxHmie1LuTSEl6e6Ws33Uet9aQH
jvekyArZEGFBeKw4zp/T99881iW3a7O3gDgiyVqDS9POp6amLe5bYrkWLgX56mwI
OGggN69Z0L+1IfvHCqt90MhdZYywtUDiM+6wt+UvWzvBKrjqQplkoUTlDesgEDcy
6CGpa/HHZAWgjj4XL6EEMmJlUF363UA+rqkD8MpFusihSrBqpOx1mswnYPUV1REB
6FmZVthEqIftaZgbVuyjl/ySN5ZSCxI8RHF2P7Q6bmr0rU/eZqAgBj69Hnbfly6W
A09+Dr6hMMksIbc5FI3xZa47pezirWIiMJWM0bCXQjUbRsv7hSUtisIgH8gTmhrh
gC4tN529HKBwCMUYLWJET8Wto/YogUArryHPkMoYFDhkmkL37iJsn9xo/F8bVfUC
Tt0vPFj3E615ukLLi83OMHB2PFev8sMbYw8b0ILmnXpkZSQkMU5lXsaJ/xS50MuX
4VXdT+51rcBTF/OnHGvi8ourx/dPCZrLZY5Z0smKt08e+5HjSPSb8iCznvlagYBu
whvUDfox1lk6cnzXa9BaAziAlZxS3fNA2sQSshEDkQyr1r5/7P247c/QkYNc/dgf
DxGKFiVu3oiED2j0YlryE1m5q1y1gUtcqW3TQu2GePrCdMcg1rft9c19m6bZekzm
vdsATuKRZ2EcEkX4ZizqnYL4E/jIV0HQF+J7mHm4lWrkwNOZbO+0nCRj1+t/FNBr
fXlOOuk46ZOKRlyEO32G2FKwcvbIgu2YwwG6w2nDAg/Su8w69oIMkK5HaDi+Xbtl
nzLNN+o8D18pnM9qQEPxqm0iIRmTjHQnTLKEQR198JvdA3fOnF8U/0IpnHPDJFg0
F8aX7XShXoGfOqHjJSF/d3WnSGfb7bPkDN/xOQ7M+qfKJdfc4fHuLFMvPrAl6buW
Dt1G1936VY/iXfM++D9NEeIJYdmeUtRAEBREcu3RKd/ktv46GlCh7CgxItT5Cs/w
m8htB4o+OBQhzZr7bjZ/T7hxXyc2N2nxZPyhA47GNYwFJYs8FHwVfU8+oKXcyO6B
Wk40jqj2vT8c1K+DisVokwsZEt+sM616OG/NoxtAbQOV9zIwnGcuza3ujWVeGMVn
0o3EH3JBIqSd1I3ubtYkwSyXecC5WY+jdvk2cODlzgmQ/FdDwfY+CbHcTxonNJCX
TufZNBJk4FZEBZhVeA3vJTRXvxhs54tMK0Kax400oLYMEH8iC4D/0uYZacP1fo1c
J/DAN2ADkt2KtRF3ZzLBDcYqFgswNrSAKawsp/xZSVyPc06sJgFnv/HsQLUSXuo5
mwXwIMiOaQ/8UNyS0M5aFbG3w+L+B/83+/GE8ERusTanLGKNQbxuRvtua/7VWI3I
tWU0RyltWTTKP/aTGNwUJCC9rS++/GLWqin+SNrLFtDb5k6AZKJponUttxtYxfl/
cjiy5JhhgFCmBfTixBlZYgvcWndtewybbAnTJu6K6WfuuY5b0gZ5OPaofBf3DQD/
oi8TkUuet7k9XzH/3ctSLwFXHRUkMCd5FqW+qJ0lneNdcQwFFB11+ymh2WM6F9f7
qeL1oHtTCXsuuqXPDqKFytYdQVtOT+mb8qTe3zeBepQFnFXmAjKaa2jHz7Omnn4c
C5SYSp+OGoQrikml7VBfGwasV9l73jHuSlnRwnI+SHK+KVh+ln6CC7pcocGZpy3I
75VZ6Ygwoxco+E4ALP/aDDzC6pt0fryoTlpVJI7cQ3vPcA2/DK1szbX0773RrtcY
0cTrP4GkeGXxHtoDMc0JbUBqyBcf1fjkUS0J59ivSciAqiM99ToRvHFsOnydgQfV
wF9bqrbb8X322A7+khfTFDgy1Xq59p+ZWkH4iMd8tr9TSWbBdWqK+26vT9WQP/1C
KzS7W8pcBjF60Ql9yeQVVQYrJHa/u41Vk7z0heib9mJ16i6GQqHNQWaJdWphDsv8
d1gRyDOazpBEWBwrrHyXUzey/bQJ9iMcibBbN4+lZfJSD2XKfDIhVd10xN+cYqYV
8xMDrkbgXHlZv+Y/X4u1xyUvJUe+VgMt3yaBmaZG4qvjvxKBmw+dori8sSQ1/2c4
Nz2umBuxHsIh79OqdDYj/2ZoosOgr4Jvpn2lNyQFyxVAGBVmXir/LXh7YlB4sHtM
NirO7QRNLmimKq47nveeGSggNrZK2V4aAKOXVGinHF0Di8IeSQvWD0KrfOzuTOLr
tpgZsPBm66/EGuRKqcMihq5WXx8LUj0KN6RcRyVrgw2ix6sq+bIvTxzQ2Lm4yxjO
elApb7MRpL3K8jbiPNc6yHuUMGdIFBNPJCsPbRIWtNISt7TO+c4F/xtOq/VepT26
cLOdbTWhYtlIXfskExWTMvkKprvr9aK9RK+5w3heFqk1aNAfu3pLRtUeEOGKO2Ns
6FURNt4aqPmSEqvDr/wdGLTXrL398z0QdGMWUxb9TgKS9cJ8wK69VxWtXIUeNLCD
2Z+cZJ8y4wEXtUTFInNkZ9wfHd1o42nTm7klrsuOc0+3nHKoru1L27qANRQlM0wB
iydeeC07tWZ8VxANC2DHAOvDXGkOtg2ZEg/Dh4Gw62k+EADTSJYSFRAxRetzozqP
/dWNYTeF3kjqc8EhKdn+aiI9DXC8QOch9cw6OlJDbmKaQ0EP1wWuMU2kIkl16NF8
mxhxFA+M8vIZCGi9cpLgmGUGVs1bPfRuefwYopUke8cGdpzEJCi1lCZSiD7wfJcY
JJ98iS1n8g2KaW0snHMsoYKKM9bgQ75/T/92I+lhwbeBu50oNN1X6cIvmqmiBIj0
PRkrQF1va7O6JfCb8qPwrFbKEuypOXioY6OYG/ll6u8/2MT+KAwt4qDD1KVqrYwW
x2MZlNpvA+htsTcWCWKHekbA68ZU1OzoAHdSfbzFTAnQqHvu01D3qrMkoekLsOYy
aII+IBPrN7YffjxLNBtQHZEd/jrd/WUq+zCmFMK117YgvHOUVLuZNPpL/ftwpfnT
G1ohDQNcs163rgunVl96cbzQUH2iSAe9ObkxJ4gsGzcwum+hI4r7jzz1bOxO8ksJ
aYbkmQDC0GcmwFz04RFFgw/xlna0fuLFRYCmPggotIYfkAVgfWnO5fmowfcsxe5K
w5SRt4XnQeuUoVsWTM5gSC4afk0mBZvjDVtpZifdrhzymKTa1Zjl2QIJmNaGE1XD
JOBXSEzlHHl5YZ+fJV8QpEAgaqU7q1gJ5DxCWoN1cCuzniStb0XYaB1h3qILfaCi
7V8r3EEaQQQZy8Z+Jj6eLKZbd6JH9cmZZOQhjMhPfcLil7sSqEn+W2t9HqermAT9
2qfueLRrb8zskMD+ghvwlHVqxyVyjYNJ4DDv/Ib91cHC6nuRV6mHtosnlvITVTae
k52w+H51Zwv5clyUUPn/JkOOyGzaWqfX0HXQTBx/ZpQn9Mk4GMY6jPkfvaTZv5D0
n1uLR9gxuTkrXRPntFbFucox7fWohI12uTcYjF3LiNous6PVAO3sBnw5KAK6cqWJ
zxBLqKhcHZ0KN91D0LQio2tjOdAUvnRi1ZTgWDUyu6eWYtW4fT8srsXgqxCBE9Sw
FhsJTNCxxJKzFDSA0Iv/VWhL/rp8FfJ5WBGyZmTEApQ6FFg/YPKqknfp3QE6evXL
uFzsP5aizcig5cXDatG5SBoMTWhc6JxSzmWLpD7atawqBnR7QnsAOG1G1+bJdHE0
DYr5VA8hHzOY9n0hhje8s4aubRscik8Wn9spcLpf5eCV7xdwRx7EzDM9Ktp52yqv
urcSq0/4DEIRW1PIYpNP71uZZ4zvoitirv9YOLIVzgjoc7isEuR6xqm4rw9OCgYE
4J5jMepRdL5LHkWqyvAu9lcAQ3B4ngZNF/8Fj6E7Anpe+xwUip+LnA2/uXmaKVKG
BiPRf1+etq8FSQsZ/MtzdSrrVkgNSud+PSwuGUEEayvDgqgpJRQw/Sbgok81ig09
SOE6EYCxDCTpO5cJeYbL6vKLhsIXSfi/ArVXOILESmh+qBkwFvNUSP2251X3L+0D
wSU3QfvB9LbSjjW8xuUKfaP58md/Yw1HgSNgAXUf7Cb4mADm+FVXccLmtwJDjGUZ
yTFf8xbg7DEvTsjz6syHVHdkoLB/w73isHGqKi2KwMr3Bhl9D70NLbOhBIzHEmXV
YjMSG/M/X0z8YI1/1Vi1prwst54vd28WSH8AbcLEmTlnIxW8zhJEeKgXdpB2cB0f
hZePXQpS75HbOxsqLmCqtBqYioxmsIuhLgDYg4iYLi15oJC80PNP3zYg75rOJIGK
89l/0q2+6l0oOcCjx0SJ4ZaB1o3ARAQgvoESKAZlheJO+90vuRgJjecxpFKuLuiY
gGMcSoB8FHNYbt6FaTpRLcvU/DYCxsg2KsuexKDsMz+dxlhKyz4dUvt/geyjPyK+
MmXrrfe4gxYg1mYKlXDB/O0u3y71cdeXqc7KI94PqCmIXzM2lX1VkBRKBh9+GHvE
QxXGySIl3V+Xr1wqtZ3v6MOuTDA8nPwuGXZBSxlQakFpH+hnMZb1OAHoygCehubb
+1McAHjegUuevznwYxD1ylJWzr7L/8QxuAvQYmdtwNf00g9y6B8kkXmP9MWM9BbL
38MgkUL+TDoLOR9NzVbieCx0ZPkq5uq7/zMXHbHCcG4FIq5+XznjnrC8MlQLL24F
CEB8+kiFKbqj502zlIwRPDV5Mh+B4FGyrGVxJIAbV9nsjhubdU7nR2Rx7fUuy19G
8KlJde9/L+unPogJnGB9f6hnVEJ3g3EVYlOtiQtYLbhYQxiTsnAK7VeERjk1sBZe
KKtumbOh/elnk7qb4xddpGftWptINR8/3WasvNcnpbmcUVSw3Lds20ICwQyu5L71
VSV241MqFKDKTlQPAVoFoSlDriqLfO9VWyR51B2NGfSeaOCfbmfIdKYD1+/X232r
TeGKNyYuZdOjNd9g8Cjaj6MM4xUk/WjL3tgxFZJkLscs4jUWEfmh9Vq0OdmeHZsy
xNMf/gpPMljoKm1PQ8MVcneh/7eI4loenqtM7NZ8/T1zgc/F+T+ROXiTCrM5vF+9
7M7g4U3tIBKbp1b9BWkvnNSDfqOB/jHeEtqeQMitnagcCjHNQzaU+P1riVMCkqQP
T3BIk3acu2bUjfup/6pp5RFSu1L3b6dBThcEDYbHSE/tdnid0TaOapT5Zwqr2G2P
Dq1QAOi9Y0oaWEi+v/hkkbn+9Bw76Y0v+LUyKaZwqUrvFHfgnrAJMWZXyJOSgj97
LSaJpYGwgm1i/gljoqE+jRF/XI9WVXpWPHT3+9dR983CZxwmKg3UGiM74aril+ly
qbKGkdTQJFNSZksn0JH12QHHjNz6ag6lQSFHohGf1EHswGVnpo9CYNuW+iIGrmQL
BUtjzNX/loKTAc0Q0dSjvM1cYH1JC3YeTY6lLrNRdSZ5s6JZaaIsqaG3S/0RK9u6
jBq1TvcNN7CfBZi2lGjzTOowxqbTkQ2ukC8tOzywMdx7aON3yfXBBMxIN6oLPiuP
JGkLHkOkisLP3fACYCpy6V7RrEotHEAqzv+j4tcbBi9uLUEx9yYCtqlAH1JrSxER
J7OD81RTOIEhFW8vWlLdsOWZnKlcRFC8D2YZPmf1iwW/a7xr04fP2KXNTYE1fzSK
TC7iwNn2o/PXT4HsrFaXCtmIELTAXrt1oVqOQPq8ePCpGMmuNexr2Tzy4SqD4ldQ
bP06k7VHdTa9V4S8YobeJ6tfOQVTaunApBF9aROvserox1OWVcBYWWRsBWhEF/Bd
DLbLlXu/9eqW6qoNZ9wJErc06dg5vy5Gtf/lt0TH4KI0IxjJaPVX/ittag/lJW+D
FCSF8QgZV3AntL2A6M62HiR57j7FsbozhhLF4F4ipL25HUFuW5L8eg/wViVQDG0z
W1Jllg9F/2fTAIQIPcxH3l3xRFtpXv6fjWxzmPe3e1IUUIpEFkCvlRKUHN8I8Ruk
FUoJOu2igzSDL/uRvoqSmZYvpH3OBjC78tCo61FedEHAuXYtEnbAjFLXHSvpPVXV
gdDIW+GUi6Fz1ilEYNgBzVnvpggNu0m60Fx28dkU26FCl5b/w4WhvNJViIhegHaM
p1s4mSbPeTkGGAy8ZMQ2fT3FZRHfwGAuS5q+h/FJsQZRv7w20MglnIEKMbL+1PYv
aHOXygafAWyf3G5BNx8OkSZCXMQvRme+x32YOoeRfSDOtB9fjMGo3WX29HkLoMRy
z1QCHYmiaYbtPF7pJRwEfQjylarDPPVcjP9Q3bLRh7fd4VxItmqC0rggscHBSECO
gv3sHcheXnhaE1DPhx2f0B966yx6WjWes1mBZ1HMEZCYL6I34WvvnnpjHZx9/T3c
4zrkrMknw1LhGr5QsAobttZbVQp4dYWqYp5B9T3WNRfFgy8aprjial+wjbHAzWip
FCpvcXU+Z8OLSUkRmUKDr8JPdFqtG9krIhTQOxv/m4tJIECEzSEj2FQtGkTVq9OA
EnH01vmohcfzKfCXAKO/G25xFBbjx9FU3VLYieAgKtUIdqxmr+UwACoEb3fKa0gO
0aLwAk+guQD5CpUXl2gjrvxtdzx9YlQrbFJgbwsSeVtIWgU4EG44BQrztWSZ+v34
yy1ba20bn5IT8Es4UBfvSsYi9LYp2hKQ/7TqrYkWj7CkeqGDrKQdOAfZY7hDCX7L
mWHYz/FUVQXD8G/0Tr38L1+UJmFw32BW+HTNCQ4wUO9IeOb8S7EZukTNvMHEDX7A
nsZKetSXj8ZnWgxL6ZZ+FAiJ+z/RO6pqsjKShn6+NqL21aSKNYN8Bw120pxfdJpT
EJgGOatUnkiddFxGPOlshvYB4Pr9Ue03a6BSs7ujeaUXKFYAfDt6vlAmVPgbh25/
dylSPq9ht+9l56b0bR7CDnFuGVnQyAFaK5+kl0akZw6zkRQuCcHM2YH13VzVKtED
dtlKKwuWKPTc23++4OQPCr3KdYGploaNCApgCKv7Ce3aIiWmBlDxAZDOdm6zj54X
MZDaotWI2iEnAcwMjAVohlhPsqjYgMEmAgqQdvVgrA5OkuApKjQuiWJkHiq81HKx
4iXfJc97b3s9i9u3WNe+vLQFb6w5Sn9BknoVIvXwt3416BPFeLlmyfUwkw3Q1I0f
+5qWl78MzZHgz/dzBTFoN7FRtrEN95snBvWDlUISE8SHL3OblD0AfAFjKrFKOjzF
Iv86uqog48Stn74Q8sGznTratc0prNTx0xtsIbKt5cFT1G+++EFzdO0RKFeRpo6b
Y2a9lhZCVXFL1FSd7VElQ5M+h8MV1DfVeZEUzYPq0FbSQeSyCw01ST70Rrk8j88m
8ON1mgjlj88xfZPK81MbkdWISbY+dj2LyxamkZEvRTEM0ixvkG3OIx39031LFl9/
RKYbdLHGaRWNKPDVn2W5zo2ucYpLv7e2PVfsYqlBjD7a8tXcXtGHkRtgUOd453yZ
rFpsMrIxOPZQD1KVe9Is+10iOqofB5+cMj5z7RbqF6AZGdPXIjtAx38DhT9h1Wua
/BJgHdjCEEZhx1NNMQdhpH7t9EfZ1ER8RXj0Py9vgC+RZ6gTb+/GzflCALBtfE9P
AVY5qw4D4fCgfGiejWKS8ApYuu2IcB6mrlQvqZH7sP5iH3QRZLWTFHsGgHuBu9hf
aY0dWOxepq8ux1maZo5Gk5Zn2sM8h5HXT1QBfAqoGLcy5pUHaZtHqjyPhsDUMsne
gqDo4vT5KtMyepKMKaULgf+opdNuhZ725Q/jI15fS1Y3Xj72MRJvN0NAhn5W1OKC
qYODSJE/QaHHZnM7mSbc2XFYvpAQeFoa4dPyd/6HF89/BfKxcp7cvXlZLx4Rnqwa
ucxB7sOuEgAlbulsrq6KWFDrxrWzXKVIWod8RG7XYpoFY1xZge1yBi+TVZ4fOVVP
yfAGeL9C/mvW5CjZfAp2F1N8D7kyeAi3jq4m+JPwtugHpHvF5S9YGOmZ5MbYe00F
dxxCU087S7qwOQlmn3VFnzqXZDff74JWTUqiHQAuQm/poAuLtEFmSVO5o/6d7WAp
IAbqmav9HaMhNiS41JO9f+hWuJe1nSkcXyW1sKWhyyJnWOwozn47k3pGHIcT9BbV
Df+ax4dn/HaBBrpFjAnBVfnqKRWMACrJiK3+uP/GFmfcwNXnr5oaBLX8ylOplqEm
Pr8RWHHZV6vwd+EI5ed7KXt30sK7FZlvev5ORk39SucXgb7kXlgV9h5sMhBZV1N7
tcdsXsRukP1wcr3mnAhYbbfF182ce3ahF6ACF8X5qaQhs6Yr639owPl/OHFCmtwC
LbkG9c439paWPdQr5MCoHEoR943XYkULv1MIMhM+1iawXs3rUl4txkU32dFBByz6
MQeHvH0CPZzY6wI/c/Mxp5vLZkjNnkLQ+2lMsiF5OvjnoJZ/gc42ZAfXk5OqkiKu
ZL0UM26KSU0dNk4l4ID/PDh0udg3QRBD2cKo+zxsJRc5v8beidU433ygPIThzQaf
KkxnVncYJcP4mbm2WGtnyR9h/pYKvsZu+pa8uQC4DRO0+dTVsBHEPoZQpiu9p+Ku
lb8mZt3hpMVPC8UBDVv6S8xzYWSCGtowZYObf5dqq1nkGpeKEs5yIQXGx2uD499j
qfoXZglBVWJmB5EG6UhGeKxm7/zhFThQ48ZItL/Gxv7jtq9ItAlRgXDvQpqgNRvi
2E/WKv1UzQEZs4x/ny5MACS8vlJXBzqY8Hb5gTkidCzYy2ZpedJJj4lZuHBKr4TP
4Wah1WBGwnQhMSZzWtvvaLAP5GmiOloLuBET5QqjdTAFEr11YAsDypZLNOCsvyPS
V5y8Jqr1RL5mbVMOpxaOPUQs+01Lq522npOSCTP1hvWJS9qFVZT2PGe6ALivqSpi
mARbjQt3D7KYjl6pL8JrqjUuyVpSKte38vHhzQmqrVAWmoAzMPxXOnXCmZR8p2rL
SBlDRzTmlmXDhsT18bCbqw/XzJiIQXFeLLBIyLWPKXqSrbsIabSvR7IRxC2iUUsT
H7/Gf/dp4cSUUK7QEIpRy0dTc854XbdlHQF55RAVFUGy+yVc5dwkp24+He3cnLvH
MDRISTzoLNJI2WIig+smJWTg1C/cA39IN1A+1FVbqr+8DC8vCmf7043/RlsBKKLP
i+1dqir4B0b+Qyc6h7Dq0OCd5U+YN06OROwRoMiLw+tqhi6F+ReiXmJUYbvEUr+z
fw0QmoqPrb9FfIfr0uIZBRoaWRWThHG/8d2yOedvgsMo4CzaR84l88j0KV1FnU7Y
6TA21ZR+7MqrEh52YRuXmwpeXaX4YoMdq9NL1JUBaRTOdA8FaL9YQ/5Yta8wWm8z
yuP39ifmBhsvIO8z0yZ5uuy+Vgb5zLGe1FJRZ9z1KGgKd8wuBnDjBFYIBMT5Ra1M
UcJVnytcLbgP5ea+nlzDOmxJy8T4oilSrHlCTJnxn6caC22KkixFTAafAbIEzL4y
UPXakwforPgE+m2iMKyAqHQX6LsLbQ+h4wGByAosIYLj42qbpxC/5MWdRR34CKRR
sbUvFm3fgL0EM+1pZiqa8ax6ZylKrmU7sLE6eeSD1jbU6MuPTl33L3sxjLNHp2qz
ESH4YyYUc37Y3eyRfN2x6QgTWf8o0piZrKM7kYajZXi7kxgnHQZf+gSluodhz2np
3RDq4bT4UAW0v+aQhp1+Cj/Ps17AiqUv97rjO2B3XT+QoxkMizh3wKbLkB8ztHgd
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
nhJr0zyz6BVsJwqdMkDdLonwl02RAm2q+4Y9PZskz5dIrJd95vt9gHcjbvxktr7W
KMMag53q1gV9awmDsmmzbiGE65Sk+kKfLgCyi4TKB2y6J6byktPZxqKxkoDCi7A3
xOelFbeUeMPgDKfFJ0tltUqcAiyAsURgo5ffTVjHiLiC9sAUJmULkjvKflCmksEh
aMaIybTuXxu3Uw+Mdfhzg8uB0wvgCMs4gTXAUL4TRoprWrdAZsK1ZyEIuOSCt7jw
WgNQxvTBybyjHYDqlz3F/IkMMpcYjahMSZHja2mXIlnKenMY1ga6MCH7zwK1CUZH
KufVyTj4WULVKhztE5HFlw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 1968 )
`pragma protect data_block
rItsLqcSZldDZmnKqTi3HzMlxpUwMfmHOogcAs12uXgHWfCo3KktaQBHnXRRPiSC
OOG5e2j3+++dgKEbjdRuHQdXN5s/F1R0x7SiObNObEiTmYxHLAfCN8vTDE68K78s
iIpNOnxjjwd/cGC+gKxJbwMeE/f6oTCJ1NdJ4TyKwL8EOCOEQAQeOHZpu8iokKV3
oCna9c4TpmBxFOOVKxAjnbYudSaYEQKO23H+3mljeQfl1Ym+spjA7HrtWPWe0caQ
kgV0h7ioxvWh5LMPNS7CuZeqo/UlicQmk0F1M5YcUe2rzKC9/cJB0QwfEZX5lU/5
hC8JsIM5KwOSCeNt13LmfxgtaAchOmlNoZ6CtEKlCL8ATNuLSM4gx3qgYoz0DXbs
S9JKzJoykU4RtxFEPbIg/fFvE6WLZfJvgaaD8XeP1p12IZ5iVrQu5+7Oo8dXj038
EAhQuJmGYa26CzppfD05P5+HOmm9eS3jFbU9npzEqwjiwJvjz/FX4NxRiPzpEmcS
XtauKsZlGajmTF1k3n8Ywi3gS9JrEIANk3CqfuP/jCpnFQQNcC0wuo8rsA/8VcaB
LYi9e3gK4uaCh2onXsGreuUxVFPI8LuS5by9bOn5qxDGcIVH0a7mYMxPqEalLsEb
o7bPkfinxECCiSyA6NBX1a+Yz7LcrHVqZa1vAIBi4ENiV+DjoJR4+RiY8rAEOg6b
3x08sjEU2oC71CINO0lcPXJYrYZqQ0OgtJBZ5BPx1Pcr3MoSvVgfgPZR3gHNupyC
bqih3G5whOVpLJgjLRozh6yyCijSfyMhsfw8a6oRU0NJD/czCAd4Vtk5zheTXeE0
XnJfdiK2VvyP0ezDcS81J8EVcKoEVVGmwkHN4CD+eO/uGDdESUrW/pNIdMwrEOQ2
FiWou9fL0ut17j3EX8BS2/sij9abZaW7vxdH8Qr8xT5qLTwMioNjHXW4PRLM0y5A
bxusVqy0OzmZyPZYT04Y9v6xn4vX3hbm7OOVeetGBY6WrrL3IYViq1zBFmvkOOfl
d97gFpsHu40ckZe9lt1C8pleuvv17OhB9xGFoeGJwAWPK8MrdpjI8NtqwcLwaiRE
/QgshS+Jt6zIpNW1n6WwTlZhLlr0X/bkqlby4KS11lsW1XkDknsl6JJGFDXgIpb+
XgcqNI6yUc+afHy9dVpRHh/TxJ6Yn0dHVHTaCeuqkY4qFv6QvPZ29wgYrne/GRGU
gY1/QHN7z7xzOdaavnuUSXgKEwaqgX3VbG7QX2ry7L7YUBssQEVRkUhd6A0osuVe
FuVyivAmKdl9y+n0rjPxlzYumooZsSWNSvfFRitlT5QyxFJ2TS44QUGrwkooPg1H
Om8VBwWHlcBDaaaQwEoDmoyvNxuJHa8DRmI9vgFjg4mdu3LXBPZ9I6YULrn59RUh
oBo8zVWU1TzfsA4+H6mfn2Gd6KAhK4V3hmlCP1100tpYN6cg+jTW3EF1F8tsLIcC
nTe2iwLeP4iaOCrs1AbN6CPAvgaZXP5Rlddy+B9nK5f8bfpFT4HaCT1dL9frM2b5
evANAmrB25tPEfmjuGofVC43dtnnEuECrsEf3wf9VCTiH+5c80lpPe8ydhs0mtXZ
2HnpUbDdI3hlp59Mi7jXz9IxY0SbFKMKMk5Ea1svWvu0qeKu1Y/UULJ+Q0fGtyvt
XoOHJf5eTfltW+mh2/NUcJdOQFq48RuhDJt62RFrVloszJ/V77sSsljjH+YktnDv
SuBe7/5I637FlkGAYCiZb//tclhXOW1IO3mTNFHdEabR6Wa6VObNb71bbjA169BA
XMuo1r3wj5DXKqzi/qOC9B23dbHsXij4OZkH6hBSPogbS8k4VQSt2W/QggLzufTI
RlXPrHq5KtZTmp1KfMO0M7XWdpe/2aWfyYXQUKFeJcwjYejd34kxhlihj4CG7Zqy
mrr1JyRVpRlOvUEmOgHcmwaKROSltzzzQHEMXQPTLehDYiHtjphaSOWikZEJ0B9I
4kkcDUE/4lilxTJk4o+AuN8S6UU5zzEOQ9ph8SUfjeUP6sJNXM4AMeQ9w3NLNKFN
hjOovnHKq1sVNdJmGuupcqDEBAmXuxbVF0VmBQggA88g51+mb8KwI5CCYc0Pwt07
36GQ85IQqDCbUPReWLy9JJ5txHVA280xbec3KuffuZA3KEaifJ2Ei72DNbGeH8LR
kAs2EasGmhs0A96a2pLdiT+2I83r5Kto4+7N/3lTPL0oY9kMAbxWLlWKt4otDiBn
RNjqsY5OORdfZfptv7ZVMBjqyLUSTCO4A6OrVGEZ+g/R/xNjjI1BNUNXxepmNtRJ
wCQZ/GQQTNbVQUAUrXpxkOY86N/800/8G4Gscn2Jognc/44t3dDJvSqSuuou8bnr
P/oDm9262IQsDF1tkl+JpR4/fFohmBXF4m6VfHT4OsfvjIaleWHECB0ndmlt92aL
P+RxrvRNbCQi3+pB9gnk73abxvOTPpBJdgGiPZ0BB7kduAaveiq+jqpWX5zuPmrk
UEte08Jdn2bZuRmGDy2TUuNd0GgVVjqQA3JOrid6s51kRnRzF24XkFcxWSMmXK2x
0Gb1NO3qW04xwL5rQVwHERRgx+oj0annkvHOQQORlBVfA8rspg7Vuu01XpECaLsa
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
JF5S1lSLH7CpaLhbW+S0navTrBgiikzsIj6arBF2MmaG20DT2a7LB5A2V9JT/9sL
S4ayIAHokwS0VsDWhYOQPEUkoO2Slb6pbfdsi5Z/Xyhs4kQKdRt5oHE2i70J+08j
hma4to5dZH4hXRdopS0BgVya4fft9aO2+pVKNa2x20X65tm3EAc1LWWORY8u9LAJ
oCoVHGtyclRGeKfFcnAvFvJysXmJglolY5fuZDnsGuqnXC03n9ao15h4MG+QSs8l
9FEL4c3fTiyMu8gAoi+sCFLpEaAKfKh5o8qNQf2R8Yk6xkbQ1auWohHRO4veolc+
iDsqcKcnOrlv0TLC7RWNzA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 53408 )
`pragma protect data_block
oMsIXYHDQMYZfYcczwu3agRop5lCq7nddjSfTU+hhPeekQaJKHLlycVOg5DtkvJA
TugP3kYDxjMeHRQ5hLgUwQcurbAhiLPPNp6++gOpyLhTbDM5/QazrDEgzZLhQJIp
wlHSpG6xe1tB/XtBUHOi3MPXngzZMQE0YsGHDwmeNYcumOqZIeXuEYF2Muxi67WR
RJz+599hqAqV++FM7AiQp990mtvFOzFyUiB+VCGkI8Va1EDS2ZUCNO3NYp2gZ6Is
pRTkDIhKiH4aDFWDYyZIgo389XUBdCY5SfDAsDsY7RsIhKG78MwR+STS8kMdkErj
L9Cmz9izTk74nOkFkQnT3QsaQuuCrp7rGT+kqM1tZlkt6EadSmTnGFnh5wQALfp9
VGF3tJwnygao/7OmB88Hzu6kffWfeHqq3hffM2+w/1rGbNCj/dmSX+QRVWp8hiqc
3rlobt9eCtGNjSlHjYrdj3WrAbC0ihDvONwNP56x17ZsJ8wazz11y6ZZr4WoxH2X
YCjYvTJ93tuV/Sf9iYpaWieJXcblsljWvlsndd5mYNOhMxBUcxruCnRh4SRRYLEZ
FUy7SEYoylgtd35/G1qqs50P9MpI0/neFJ2w8+WeenKhijmqtWPNEolBT+lMn9JY
FnE0lkacu/2tZOFuhC1b+woUDzg2TbNSE5zcsISGWtQTDO7QIonjgLQ4N2swSfbF
o112Fnlmv+Ea9UYL4DYYBxWWVmeP8KbNmgK/4VHEtxaryVK6WaGQRvp0WVIDCu7J
EnVaqG38Ev8HBin6Gx17VmxGNijhdrbc/sz3Orhpql7Q6af2dcPxTVP5jr4aRt88
4avtdljMxXbh2FIoRFmnvQxUZY+lfEulpMqbm9poHlJ86QXUN9yFONxEyE/n7+fN
+qcKU+xFLZ17m5KK3H2jHAehCgIb3Qp0GYmKcNhPfe2o6YRb7SXYNhdEQNIopIue
zMhyxYsYDdnDedKYD/bluDsqfPjdU3mT7dol/r6k+gGC1JlHjE4V2kvqDoorftBt
09T0lNWlaCmCYTlH9JX45d2hwE2d+cbtZxUizc7fxq+u2EGHBcboeWayeaG/2TVo
yxFJtnSDCiLi8Wwo7nwUHAPXqkC3pOHr34r/sBs0AMP+0Qk5KDnaaYXL/UlgbhQS
mCzneuKaDb9WT0EbKZCxD/6Q37081tzN1bPmZYOmJeO6bYxIZ2lSXIFqK6bhl9HF
mPzDliWiQJsn63gOuQwYpLW9HAKbzTQwJIr10ogXoH00HZ15THcwZuFahabgsgJb
5g7IcOrH77bLJjftaeEuYGGRqRltkDTDBsZNupdAX07jpt4ZnYH7cZzHu0DLiifp
hPhNTHRZ8n7CWsptnuL2y62DtIGk2c4LnQsoSa5OfZ9d3qJB/AgHdeZNEtCgncuh
pLJao1TrLT1JJGKb6PxjGghItlUcqU8GSynUBMdp4Y+M87EvvvMSys8J/tXdePO9
k6ymm4C6V8molk8o0JhcYXr+Cny20C0ZrG5YiNazj7uEBiG78P6GpsGkWgh6JP4u
yhh0v/+UBjv4jxQYQ5HLMblrNmcqvtXJ0xhmZowTAL+b1Wj9VWrgZq4DjMhX4MdG
yHqbjnWbZIkOlljDaObKAIy1d5AyUUsetfUxZ/5hkh4kvtW1R2hGqCZuKleUYooc
qbmlcTP1LJXXvfxFVxBhXJ7JE5Nf1HtGbl+ukPTDsCvSqwJVMdBfPsFBM3RQPHN8
gby8zxNnetnl4m0OnVFF+3ScTsqEljSDuwm6JfiqgHsE8qKW0XiRMuP70KIsabuz
35HtKbPD1wiA4y+xcmHjHTjaVU8N55FobkWxle6EWD56oyUJHQecrypHFogoZkQr
cTmeVLUICIXoEyArSQZ+HBv7JYFcUa/SEpOMBeFELeW52v+TKYjWLm3Ycr8qGdQc
WqGJE+Lmm5+6FXsRZZF1w/leM2KQN2igFgNRwIVO5ncIHPUF3CJdAsIV4o3k66aH
az60lwhVGKMGIyI4KNhYrLMhGExg0iK1roTOcGQnkVx8qR5cqrpv7AuRo1H07Kxv
gnH4GU1iM2BfKTDTLsV3avabGTDybJrZ0LOt+Y0MDlcvuP2UoIGFLSl4xGk2Xgp5
nkoat+oZ24Gr862sa4dYT+kklh3R4vB4YxM7sLJs5fh3WqJ8mRjzWAtbgVDCKND2
CBYKE26HlAaaxQpQQOFWA3NfTX9/pVzLlUKEnA9q5RGrLQuQaFjFjzElqaIUlEuQ
4U+H5RzKv2iFSRZOjfIjFTMea9Xz+iXt4G9m6ekj9SFGeNIFiLihj8vQ29kbZ94G
ujiy523bfNLJG120JSgTzqDKMs4Ie88x39SKHdm6ZkSkWMfjW5opdiOKExxFeoYR
Y4Kl3v6mC9eJo2N4f5a+BbUYcHs6zpcoQQOGEpVToXvfptvoGSlSjECadzfQDpyn
DLV677dZObO5Ire9+DzV2MWYXn0jNPFNap0xKn/yw+trBLOSnxZXBWvVenYgE/lq
ZggxYLGyIW1zBkSkvpc97sUrsl4F6eOyNQbqG2fG7DBOAslEygf6wPs/PIyYWaU5
di0gOG5POzIPFclFd7W/8Bf3xaZPRrN/422MdLVDjvirzonpaGzB82mUZaUpKVir
Ahpx8rjU3G+K4m7yR3JGNYqqMx78Nq4KdGTg0FGPPokRUsZKFDgvicz4lTZSxrYd
h3dfF4XT4iSZojQa0qjQl88EWZO/v6Fcr8ToV3UHVgiTHTgg/C07LLm8W5TT7NRD
QJfFL37f/Bla3zq5GBTg2Vzf7ftU6LGceeWkjMK6kXsJ5n4Z+v4Td3zsmD8mFE9o
dh6cZAQDqjZnBePwdAtsa4YaLwW+FHHIEpiFfXfx6kRyilxX1yvqM6S81VygMIry
A2d8wliNCW25DB8KFdW3kljD1aJ2xnzevdz/67X5Mq/S0FNUhSKfyjyAL8NqKoGB
yr/YkGqAEhyTeEVdptFnJv/P/Yy9cuew4tugB6q6kzsaK84fBtXRHzOkZKGq3F5p
SqmRCm4WOSmH/BUErnNM3Ci1QSMvCg5h5xhTYRSnVNd41mtUvQoNmE4be6Y0oLBd
2q3jhQ3959RUO6St6zXkM1AEwp4PUz5jMhB/qSuUNXhwl/0aC9NONZ4l09jxmcJr
M6Az4qUmjqe5LRY4CLxPNt3B674dsDNHbAgz11TeoP+xvGnYNaeHsgGUKUyEd9En
GxghKY/XvVfIIRdI+YTrXAyEYnCjmY4++GFemFIBoQOoocKlnQHgF50/Xnr8bczw
hpNs1ebn0PFWhgtkCiP+UVCMg6h4cAO/HQrFRym1n6S6xQmQLVZBstDmqf84Yl5k
+k0SLbtsWufzX98oleOYASMfnawxs1FxGE8dm96WhtQ/VDVryWYzQDJD13X4O2Er
emo+vlKULoZFwfkn99z82I82eLPyoa6WmMyqIlngOvco0mF3nC30ewRVBlD9L4yl
0HgSYCgt4iV6fMsgrg0yIYJ0zLbdPGX+upWlOE58dnqOmxa9T0RYB0/6oFwBra8d
IoKwlcyfwRkjCJ/C2mrApI+AmYF1brww0fvfb6QY2uu7Dh/cQUYQGDz/vGUXOhr4
8SLwkBsmliysOsXbiB+fEloTAiUF0hYdYt8aOLAooMuGn7EehsjxE+RlMM65eYUK
fnKBB81DdkpE5KikWSrobXFeU8xKEK6GYnywhDHh74hii+RX5lbEy4hScEADrt6G
fvPTLPZBj+x0qIxr3oaPmsT+Ax6eMV6rdb4+sRPb/E+5pgPDhLodg8kqNxw3rtJD
FVr3kk0l/8q+82hwlHxpyWgVsxMEOtRILHQ2dGTq+IbpRxm/FkyVDZaoSjrBVlfi
LAfX3kLT049QW53y3eS4wDV2UCet2PxYZ1rHclPhmLc4vWJXVHFk00KZToq4Llzi
rS9yblrf4e63Y+4Ws5sWMFp4PYbxyL7k5gpoeyZVMxvATxxHe5uh0vuAUXgN30X7
r8/mmmEiFM94243TxeWfBvgTgAd07LUn3+yDqdKEAyFj4MpXXGgJLMxdrL6vr//w
tyAljg5adAPJEE9T6o5Qf4qa0sbylgTM/izO1KeWPV6RFUWff+pUwLxNxB/p3slP
SDynIhls4rcwNtf8iC8wG7Dg3Vn28SI7UAu7q/+6FKAlxfAKz4e6IBCyldRWakjm
VMF1LXb/NSdkUV2baf8CEpPwuz+NGG/Tv9QlavykgndLGZk1Zs/yKVBS6oNzXbpS
7uesc1EON1LKVxmXRRpMT8E98T9amFOOe3neY3ZWw211FRGUP2kE+dOFuXXeFLZm
leg1Eh7MaBrpCw8ugKMGtIJRnvWH9GR7BFJYPpWJAz74/6HCmnUqPR45mBFR0Hj0
1nSxR8E7N9N7XZwcvJ4gNVCr4r+K1VqUhlDE8ZZx60WX750Y6jw7/SKzQWWu6e8s
r+oY8+LxB0lHyiRGJ9gSYveUuU39EyjIQLr+6yxoJjPZ74CF/cNK840YnGc5rZUf
VSHxujwWp9Qx2qeAaTEoZ2WsCpgMlV7vwlbizalirPW6cp7eMwCpwrIxrCuL9OdU
2j3NmNuGcPGTXOk+ekmRLJaeLivkVOZZxWo4gZseArZAzvxwi2pCl5NQn4GOjEZd
Eq7Q6q+nkxdHcqo4Nb02U/mk6Lk1UaoLbiNeJ+5ow4FoOZnbLyj/vQvxnfBXwAp8
iAVLKJ+Sg9qllbaF7FxQXkfL86r/IbXwR7VP+dji+EA0B1ZXh/xNkkiI/5ksSTvP
QAHSxsnDD4px7B1oNQ4p/y2MD8nDV0H5a+piVe9ec8rrOMAudocd5TBkzQAfL4Fi
TE8pw3na1WXmgftPNmKHtlRtQYikrdkd/RPPf+V3tbj36w9Hb9Ch17rpyt8WxotT
yNysrplqVZT6W08tsrCNR305CjRSZoP5hC5/eVsdztsw23JanKWfi5+xM6pH6EYB
My0eXeurtA0UjXJDvmolPpDnkFcLeF5F0SATrYoRpUZlp4TN4D+/Om7lQFV0YMQS
e6npnssINRwTbBkoIsQUWTPhAWs/KBNBwKKMq3fMajPrXGMwxq47jDz/s0+gz5fo
WoaIgxLCtLhpo0KoHVNxNDNuCrCVdz/RO+s7VOaQyN6cR5vNFZYapTnPdSs3AbWn
oOp+QBp7kJbfLsO3jMpIREIe/XpuALKvdUsHX12YayBzhszo93Hjgz8QnG3OIvLL
uZ3VbYIg3T6JogXGZ81MIADXdvDYOrnnqVmETLNN0ELbDDRC7/QGmFKTtNJ5uA7Y
p0i06mX/xKlhIaFmb6VnkpJGKHlTpU1lOJKAeBFBEzvbuvlJsL3pKWwI6ONoKumz
tjwzdM8ss+tR7zRf/Tfr8cO4jwetnvgMqCH19JuvqrIoTADJF03arHZ0J/AJFOpY
d/twna1nW6/Pnr3EdFzyoUVZYThF8x/q+ZL6aiUzVGNah2Livau80Quukg92TEuH
EtpLDBgDjP4XZEVhC4y2WL/AJRBD4FHEX5AFI7LT09VLHQ8iXcw7tVY+VmF1/D1i
XgUzShw93EBhC42/Z3CWuU1tpJ2h7T9mocnd7TohKoW3rcq6vZu/hKqnUPpIPG6k
QqqLyFJK6lSIRP82yP38pp2D2yuVRrvO8DEaCfz+/Vxcxx58upUi3hK5ZKHYXt0m
cNdXzRJV+SGLlP74iiSUPlNLOiZAoO4xIcuueougsyBeWDHi0Y3oVKFp+Tt47SuC
/+xJknm//jGIHrQRJ0I/BxP3mq/l2+3aIDjySdozfcoUU204KufVOBYOlVm+HoUG
Yj1Z3BpgUOlpL+FA6QLrfPetkuVlkCYtJz80477sK87EsBscjsBhvPWXuRueeZ7k
mcUBjsrDNr6hlBvCvb8Nw2kxvZ5R4f8S4NPSbLjLi58rCnG1SRVZdswiT/ZCOBSW
xP3d5Sk/dDqFEN6Gb6Ur46eEL8KFsyuOsGFxBIkwt+F/IMCxIBhViSYHj2wCVOkZ
4EI86T3V6PEZG4ICPeF1DnRfQsza3swJj/7BTBMegXphrDW/xHSar7NiPijqsidq
01FamEJNuGNEte9Q6SfkUcUow8wyAelZ45DsVkTXWOTsTjuiTswJ5CPILpYt0QYX
RmIQjXmfdIWNurGH5/bfHYW91vloTD99w4jvfrXPWA7TwBqgtq2Xk3YmY4GnE1/M
98HvwiEqj0xVgJl+Va4dskk+CEiiwYloWb+SoyDwp1Mf6YDGYbo7+1nh1J3647a1
e2M+5/zHRYPIFSnKyfhMGkXeCdK2wMyRP1uvermlkS+f0VM0J8cNHANt4McPzeKb
feCsgUFQMfQ3PVpYtXT+DDjK9VMmQn81yNjyKYyqa3VvmNNBlIJqFjZspUcXLW/I
NfbCJZz1JuIARJ6m8233hJ7+gq5A7SF/spn3m+f2comJPYXCYvyd/iQr1hhm+900
r6x0OGX9/D1/8cOH2uP6pjhenkqriioPdh0c2/Zxp5upUi+ny5dRFJ/qLeOXMOln
ynRglW2GNSYMW8OodtnYLQ6WYxUCysrr0UjCQFyQQa6IDa36nG2EkgXmENXKsNQK
LE4jjTQ97OZdUnAMEJJ//67wbFlKevzuR8HiLGIQoP5DLsNf1sbKggLS7AKb5JEb
112f4jB8vyogWrc7PGXwQjJoz2x2LYvPJTbvsR2Qn96EHKOmsAyiM8Tw2B7BUWEZ
1PGKvXEfVwiwBHpfih6Rw0fVzMia5u0Z7godW000Appd+Fs9B/ntdN4RCc/ZcwFK
UKQ0lGa6fwbv5gsVljoA95Z+KQPZeFZAtlNHYtOkjjEfVNId0RS6/WfWoTpOf0Sl
KTss+C3FFonlqcC9EgZF/ur+qHlKjTo/81G8cOdOTZR91M66+Xn24YyN5Bp6+OcK
25YekPd0++LJphLnp5iV+3K3dXSpH0VHNuoQ16UjgylT2OFE2uoKeceKAlEGkZaf
YhgssS01MCLbwY22q8c8ajWeBevyI2kzS7Paf3xf8yF7Fz0bWcjDmXmn8eGbx1+n
jnkkdWZM29jqCEkhQlf/EgIQb9SbIkYpvyBYJAcwXlaH64enm98QJ+xoxdJu8mIV
DMYp6rclp+oD5qKhg0FijcOUtU7qIvG3uIOCbJo5xhnYB/Ug0GShJmozxaPGpAY1
tVr3qHpcz4X2VPfaWsXwy8cOVusr3JeJ626PDjhBYwzz+UXkSMPUwJnTcy+EZV57
9c2ayHZSmin9yEnNoHNSnyJN2dD67PBu3RDgdbOrsydrZuBUrE0i7qfKNDHWYBb1
tuR9i8hMUir06DmBLouwp/73CKaWvcm8gdvlxYr1QHJkkc0BiQwqmCBRk2QDVfsP
7QqLKtvFOvR/UjWTpyLEn47CQyo+EgHVjXVVqLlvg9Sqq8cJ3cx784U4/dxrYRy/
VjuZjrMtLRKdbpieFL8mlZJpMPp9LD3Z/m/CR7ZdHySidyXpKhxdm1GBgffX02HN
fpaSqEU2tcFvGCtJ9VvyWbv8q5w407lHvKqTMSpODwY/KEjJd8qcX5ftLHZN56/h
oACMc5hGIV3DlaZA9Dvdk9cW94X3ms2rgYei68V7LUHRzYE3B78jb0ugGjSXB1Mh
geHb+XrqfTB34B65DinjN6KZDWrbhmcdC4dQoS9WHoqhGO6LhDhXI96tuadZkS5c
i0TZMYxHUnIhEST2c4RoN55cmpP/ZAPhLZ/psrSq6ectylVHwmr0+p7iW7ezKlIg
z4URdhSxz3TgYx0zV6kKUizOsva7AdCscvKzvYv3SingKXRQFJ/ZeFQbqML9WFKy
ahbcnNTD2HFW04cwBVExa1TBqNGNTKY3ppuXXqSDJ766gccYQM61YdhnA8ETgTRb
fPHl/D/PANAyJsyzZly78lijbVStAYYsU+870W4eesimbejlvYyr42I5RyyQ7B3m
M/ty5SnYfH24N0+R0XXnfzk+y/6YhETooJvMioXEhBLok8Q684EqWHTD/2IW5GvL
cfr5hZdH7NYErQFx0TSiJ1XjMM5CBwuTGQNdjzo+vl7xv58HH3I3IZyZV/EtoVWW
xRu4CKfGhU8JktNkityefaa08GsXlFzyWypL4MGFiN715Lk0LYCo9LJjrltpnUtB
8Me5ZRp1ihATSjU856OKlUAHq00zMiC4o4Z141Tvgo2JhxxSVZ97+tvmQr4tgNM7
47MZPhuVUnZhVQfBdPMuDRjy3EpxQeXjgQPdwra4U5fFgwQGrrQ9ft8rLoncknBO
tfpIZJAadehDQgEZNKsKZRAvp2N7mI7T0+xCpUTEArIRryFI6o4se3phpV7gSuiK
YDo0rH8R3kM2ubXIJlLOzU7Z/tKZYMV+mxSPwUxFrOa6SQXvhzOhkCGaeGHPs3Mt
Z/9Ifl4CZKyUolXGiWUAeFulqE3XZL9dFwxUCRzhFCGyL1XzkPNqHnPhzl9agzHY
kJ69S3XUTjDzCV+Uasg52GqAb/ADfUHsQF4NgwqTTF+IL+aynljQ/hU/xUFtBPP0
gXAhonjTFyvW/aphYCgnk9Vl0CerFU7vwzImBJVz/vCZz1UhCLiWtNsdI3nuriak
3rnPtu7wj8FK865Lw3BSL2mD4r4DGmlneK8TIu+spQxkjd5D5HsuMCrnaMGDZViQ
q68xcJAKUesyy/BqeK39wboUDL/iw+CO45ENgzCZHWuT5MHLMQLU+l2AXGKEUj1a
T5p1MWkFemEqeOhCr9OK+AYSUGLww7AihU8hqyOxJYf2/J054YF3jn7/MoK1kpHa
tsJUWRPQTNuhW8TG/MPwoTSpslVG665NwQC/kthhdEMv16IlT2C99q6aDs6Si03o
GuXjNX8T3m4TJUd4yII+RZX9hdcZpGmyE8mYBZxBP0A0QG9668SkyQFIDGLI3cIi
hKawEsjI6NL3JdjjS6OHcM5E39/akTUaAn8E4qBsu68SMOoAR8AvNIkLWC7z7Zle
Iqw3pQYRcmg/xV29rTPCMp2MQIfH659EYwWcjqoymOdN7lfXVq+f9ODu79hUCadt
gQRzcspYci+pwCajmBA8mtY23Xei9pzReLM0O/0PL9OZMbyD/5Nn3XIZQJe3W1cZ
53s5CM261uL3bvleHknWIKp91FdDjg/q0kRN+HNW/ye7SZdwL6YJ4zNfJEvg4SRF
NTlDHkBj/e7i/HOkiEiE9w+5NGIpZfbr8/nXsF4axchL/E16s1m01ntkym+xWk4l
yjKCX1JDuQQhXlJCEVqKt6d120qf5vSXUu2AJUOKi3KylB7srlQuKfhOIoX9RFd/
E5+Dm6Z4cdwCx2ak5APzFmjRiaAG6QGE8ibLHuD4jNru4vYjv6UK0CSLqKeDUGd9
YaDv7tFgEOuguNFCHtBksSAnFqaOIZzhvlQY5yjSMN1t0RdPF8IdJRAFbSxFObp0
5XiyiaP3wp6SJhgqiqvUh+vdCIzyhtNU8u4Qu3XW8+iO4/x/l5SZGAJ64mEXXVSL
ucIPSswUmrMProY0kpmhsTc2poJ5bALi47YAFPRZ9r6HTxkRSEcHFezZirSXr0PD
WW3Q3rFnFENv53pwnaZc5uanQlAlxh9QKD5EvrARoqws+cznFO9DUNj2EO7T29Nv
lq8XNDy6dFNfe/KSCWtPdE9w1QZvdr7VPH9BMRJ4yai3YPjiBZVSwPt0CEQrzS+y
dJDEsqM8d4vjPuc0I546zfRf9WrH+RdZDrz6RFDih7Qksd9bvzUf3lmO9qJNXh5N
V2ZBlJtVnZm+l3FstBHXcOfhOJWDXVYpsxGy2ZGODb9gQ7Zcd8/zL8hcIRRptaOx
fy9lTamLRG1RkJx67q4x08pK6SRssCUsgk14KCwGDJPPj/EaDEJfxEtOpcZV8xG0
8m/jOyeFgtvxAUKOJfcg/Hsf2a6I3y9sPCGTLxf0yTNVutNF4T+o0XJQ5VvYxXlq
mai1hpHI87sTsVgCRRIIWDwolwIOT2qzniyc+1mmJv+l8WVg5Be2lXOJZPreZ7rD
M1qNN1M969fB+AA7XtUXOtmqKYccw2CRq1syCCeBZPvD4bh7Vey6OgJ/F7LTZvo9
dWM/MaRkC+GEYoS71Z+EBPjvdfCE0bpLnVxDjogAV5O1MFwQzudowmetJM+Ttjf5
HtMkUyWyBH7eXDO8fINXUsNqtA2y9d3ziGi574duIRdGxZyz+pm9A1kCJcT2IbSR
DdofJ9XsRqQPu9uy1nYrNNyE08DfwbafJaYI4DuHBCnV0FTNqptzQEYP5ViJBDT4
I02RgXCzqaPC2UZqlETbtvgD+DIRlTMRprfrg5+YqGmI0xOuuC4KgmXoX0yjfLpd
qto3xFPHDFBzUKyMMcxU7RaNtwGS/nNX978BcvAJR0SP65B588HcGloBgygV8C/j
C/Uoyv9s5uxLzU8dRv58LQHsiX7uSlTb7OcBP9d1JeFN7KZTfak3VH+sVvPZa/2Z
8IGiCWQaX7cJlQk6LusRNtU0mi8nu9k4h5zHknMl+/fqXrbZPHSoHARGatQJqFYf
3aCbsoDerTH+DUf4ueOV2uFtlvFifa1ZjrLYZfgJ45FZSZukNDQGyve3FFOOK+rs
KsrbDoXE8v7SwylD5IyqfzEj9Nkczlvbi06R+eeyc9H+UnbPpq/h0Q5ZyW2MyhIO
1Rn6EfIPUSQG/fHNab056dJ/v3HtFkNGAD96NZnFyPZc2Gn267OnNAYUL4irSGUK
zuaDP/a5qEBATL1JDXz/v9XPm7mGITW+OfoEA109n0dIUJHX/rtYP3/qo9mEz026
j5IbFLZd2nrONBlKouHVZVzp8FTHPB99GSERIQzuHUiA+XSHZ7Sv6ls694w4fSu6
wVZwoJPEJL77e6d6vctn7hRd41/6dTlI/RHEFlCzbGMF5gn2QLr40+9HHreBKvXx
z+XNCPwSEgihBca6EV+ZEy89A2Of6q++lwEKiNMU8CEZt25JAysf8kCVId+iubL9
SLMzBa2wv91cZUMTl6Hb3SfJqz8br3F1JOVcu76gmGyWbB3AQRBCLUibDxgw1QdL
3ShnFuLUNrABUvLhWhhZSFR3ehtB+FynuMs5rnFlGjilrho8Ym6Rck/Jy62y2kvi
7D7eA84iqOTgi1OFXqZhLKtSYs3HIgZJatFAMdn4XGQrvO+4Dc4KsaW1MxigwXVf
0rA75lE98NxuuB2eMMGc7PNuqCBtHZc2ZuD0id2CDscxAFZfuZVFSLtuaX5uIVZi
u0FT3gJfjEM2qW5fLqcOiizhpsrzALShkM11UOXK8WoSyZ/9AUvHtanH8snqh0Yq
7jrYF8CvYuAvIqBPgqbWbZXK6cd3THtC4Q2pVqG4QyYEKQhHWU9HTbGtkGjgDf8D
8K7l/ub+ZDUm/KcGpWfSwI7bhj5XbnHu9t7hiK2mFkcVzdEtBHwdNMXLe1My2AJJ
cHcEnEd35fg65u0PW0SpHIFQJJIS+zXThSaa9E0vAyVWI52F3is3kOlDgbzA06sA
uSn6VFYVpztROPVpvvXZUq7JbV3oFRxbi1bzDdy6eOzYkX5J+gAL7n6Kh0P2NtAV
NHKh6IBLPU6WVmhIXnpzKqc2/6DI2149Y/v8++7HUFdgKilqnYz1+nPCA+FyWlrc
H0fM/dgPeLWwsedhxT75QBY4RCaiDu3Tfv3KlA1wj5rgEoeUb3ruQAjoTEAgwzB/
dh6qu2eBhc74gTZoYuttNAVtykKk6rehyIbvUOa4NX5/pMTZukuMlCJNpMAlMRxW
d4wCFiK6agxiNYIKn+W1egTg5ANG8PEN6tOCcdQCNXR01oBwZWEIQiQ0fj8F2DH5
fp2gw0fUFGEflFe7gaxr25M14xipmOSYaqWgVcm1Q2mr8Fwcc23Wdd6L7THu7x5A
IaADFcioajNsuGA5h2g6V/rByGB3aYoRUTA73IqeQn3rZu9+Q6RDKaO5xBPzjdke
mNhXYKvu1EiMSUgwojVda5bxFGkh0UVvQuC51jh5h9eFAZEk445srmy4R3ID/3DW
CoezoZh5+rzfiFXa0LblHkzVqrEo71wEZd4qiMGbzp0hVHMzZGaWE6Kno0Z/ivMt
zMknu80IQrYZm9bykTRoA9tiEBqor2oKGkxz1bQl/7BIsavm5RxdLgeI0uJ6pkQc
CQKHs1cPdXmGj9DKit1Mu/pX/1WClNXHKx/awIg1aJlvqgxcqrVFdHLW0qC0/loE
JRJgNryBOiprCVF+veIPP/vc/QbVvXCUirytHgUZWvBJ2nePUi2EO/tdf0An9pVh
Hckpzhzd+g7j+ymcx6eFeWQtzwVgmumI3ni5lhgnssa7Nj00P2o2/d7KM0La8yvz
wLAWzH0qHzii1tWwHG89Kj8IngbCd9l/cJh22zJg6rpAOEPV4CE1O14FvhpdZYqE
mONuF67cQEUqMzLtKh97xffUGQ7bpqB326usbd+MB3H41EW9ciQO+Xgf0Sni9soG
RwF8B2sim305+KI6p62tyRnkb1qI95QQsjgFrd77VqkLPEnVtGPi3+wFcRnc7VNT
P9k0tXJEmA4jVGYipr+oPMBMeCy0IZj6NwbYqMAixAbvnLq8fS/JVcUZdRrMG1eM
l2u9nTFBnsXYe9DYCdewUQZv1fp7ak6BlMD/MQQJnO+mME0+K93H+vkoMPi3ko8u
hu3W2Pu/pZ2qlXI14uKO8MFIm6fkDAjdAAhK/hFDBFVHx8YJxDWleHD4cBkQPEGX
pPAqXrJjn1zL0cyZ96BEwqueePOYih4JJ8h+FuEqQlp9WfWsj4cw/KdPhdSoPXTR
KJrKXV5lTjCfwYpTkh11VzPFnxK/CwD1pBW4ecs61X6KkXiVWkrL1TJWs67F/uWB
ajkFDSjnfoUihmrr4pArhSAFL3JVPjpRByqLz+Zu69amBSmyfDEmVQcvjtqbC+Qw
BQa6rz8xB+rmM41N6vl1jc2pr/Yr9reoFJrDxRXWWU830beJYQxt5/njezapVYOG
wVbW5y2QEwbTGVJHY3qswuos0oHegvuXOaynIqHFoecSQyV7i+KvV24a/2O9bD7O
JZmiV8jaZvEaOTFFt/4GjVdQ8pKWOy8vklcBJVroGctD5yq+vL+xjtbr1mzmvhwT
nltxtbgpqJwIpagvOcSot2/kY9NAmhDqaTpvpqiS/dGsgprQFsiIKH21SL/usB/Q
bBKxwUAYT/bHeNVY6rlZoP09X1hEQDKf1uKb1gPGASLBFrx29o9SU1/mfjuqWEmc
cFwYUzE/LYERtCRgX3n9xxSVrQbNVFROjE+OgauwvxUskCABVMarxEcw50eLHA49
HwlhTqY9AsaDys1kezWzrGiGp9WMp6tlk5l1nsVNO+CnWmCH4KatnhB3YG0PhfPB
sYPJdOhb5LFTZBeCiQUu1xV95ID1QoXy00KMvqRVIE5oTX0PZM4PinZehZQ5JN4a
kfXhUJPmgekQeYYrbXVxJZKnXTEAfn+C9KOfrKXaIIqETVwcZQDbKMzclTikxcmT
yzhczBHpb/RsVOarCAbgQTPDTPQ7kQNAZgc3ix1Qn8ZTJDu1dSma1OdIvVC2TiQ0
cvVsa7Kfn2KPzZBLv4gcVG2ba0W7oKyVi8zJrYZXiOJ6AQhn7V6KaXeA5roHf/ld
9xUF3DQLPWw8qrIAdllJUhCXuRTZm317bdY/Y9yxuw6YGaoKSCEcEy+axjMxUP/h
SAhOrOXRTCEyJQG4krjRYox/+xOClE4hiq68Uwo+GlSyuAEvRG31FdjHdNG7ICh0
lcIXOr+lt7zSPtmO7q/j0LAeOfY5sg+Wn0KocNcCDeQG41WxrJIe0x+Yz7eFzLn+
5pG2fEORiiuICShvQrUwtwk5gNrYLlP6sEzctFe3sLxgE598dPPVMvR2brf+MoVw
GP2Q116cKNxZDvNFs6KbJRrYyOC5dxpzDwRghJdQVO7f8T4o57VwUtbs68sMas0g
wy6ymTkwMblouXJQdadv+k4p0OszLBnUy5irYBspTUdZlsEcbn+U2O3Z1UN3nS4N
AM3dAzDH1vya2XUN9Q+HtUYhaguULun5+4kosv4b0bUE4vbEX4xY7Rw4bQPzdGNf
uVQ6vE8QQ9YU6jOUq+o9yfsHPrE/EtARuhX1Aq1+fRkhs2nFs5e8XK0l7/l+8oPh
fNlSCKcNz0UzpYu8bOMDz7njzOlFHjxUnruAgqHzythkhFHW9HjfTfnmSIs0PFCO
xGKoNpuEI6+lB5zciXHE+hCu1Dhz8hhAi0jghr+Yyl1M6etPZjA6K82fWifazkXX
kDsgkX7mauiTodhWaGCvW7OuviP0r0g9lQtJcxmtqnRl/cm42eRh2rddfrc+3FVk
K3N0ulLbunZT1ykds4iTY48YzQGUCi/1DlFSRHul660JKyDH75HCikL+vZ/rlTGj
qYzkeePll4DPn9lHIeXvWjVMPyCgB2w4mp9OGk8dW8k+TmMd3hk9QTlEmudYp5Zd
YglG4zJYzzHcreBNwrtF3tTjbMq5xWEg1diTbUBajpv65JCHHZfrViegNDkliocI
RDUXa09CR2JJAiBvRr47KTrgtnkT93Qb/Q4LVunVJI7zCq6jWJEGmp9ePsli/I9N
g/GaO/wVwZUrPe2t+Q/uqSeAMn9ff70GaxrRcJOy5Hol6VxGO1PzrlrzbHnGcvJF
SfMJ5Ou5sc4o0SAODNkA9fvTnd+lpuBkF8WxmFHwubzC9+n7+gXpkt1GU8eAYEFp
4lGzNoqAKpEoOJtNzdW/+kMCYt6Xs+J5NWrC1wI4+bTs/zn93rGqae9Fs2jvkTZD
rE9vwcU0Uv2YkDDkabxq5jqhHcHCI0LjfUTzIy5ZJSPC7j9T6i9NlMLxRy9GcJMc
4PJTtxSLpEkkxcpLTihZh12B6+yCAcInzl2gLowvEPHD0JS1H1plYuxpyvwPPgaG
vQxHpY6bwmFO+z6U9t1ZAKEoh0vzHmShuFNS+K1u1fVrw9M/9ivNqRl250PaSTKw
BlQG9A8CZwIOEJVV92LVM3Pa7/Azl3+NyEQadw7JtWZ8eMN8fluOiq4UrgBpiDlG
J/53unG2XHzwDwbutXtOiQNJoCO3Ux1EsIPpxfx1pgJLRZme5zE+Aq7V7fg/MaUb
IU5MCq73OwngJXD0GBoQNpopNuNF0UfvFGKkRSCz8HV882Xkho82tnN3qOwBANWz
KyysyvV2EZaGinjIAGL+uvSo26AYa5GlmfDCpxZbQOYBnjzm+mGJOjoin+i8YoSf
fRCFPlLD/Aa4znYIp7FmyDSu24ELK8+83s2KWBeXNY+Zd1EpC8520SKKSAeJg4pl
zpK42h50OHgnQ40/RV4lnTcIrYhLQOxTBVHzcxNsPYpil68q2TngQxM6Jh72SFR9
lBF4iwYTtYszLItDZ2MwKgseCeWAcLdfbuk6JMPVSlhvugjy5mEBgov5dw9NCswK
OHnLgaGMpUwJ0Wi4OVNwYrAIF7uFZdizpHKX7ifLaawyKYJSA3zNHQlH7zO+3UZJ
wbp88Hfoa0ZOoZwjvDNfM00+a5sNJId0nZgVxQPyF5iYAW2CTj2naHlQ7go/hKoT
+la/7lJbIFFSZyo10NJTWKtMZiPtlwuGUUHSybPMYq9DT3r4cif6QJhAHB6YXau1
/ROp6KPmmk683I89mMat/+UnoukA2ojPl1q7UppB/BUfer++VSpIqYkLi4DjT0az
2EQWhdxM519tDzwJt37KWBpB9eJaGW/KoOrfOlJQDE2ERGGOXQwlQBTCPj9CcAoa
l5lt1VOZxuZq92LRoX6cs54wWo2Ok/1hPQ2tW0k74/L8xu9kRiURYMHzjZcDi9Xk
n6Bmjg/Byz2DtWIoyE+OHluoahp/XsPEEsux1mT26Ww0B+G4N6+WLJa+5NuqQxWc
XGMC7XFs3rm6GspKWy0ZRedHzr0YEX/QptBd2/a2pSA8bgnv3zVVfr27bXN2YWWY
rDhaOeCvZtAwfWVD9SkqsCeh/vSUhrEVKAcgHH/SqerkrV0nyV3kgckyjjNeBxed
lrP5vPHApU/uzJaZ1aEjHuLLKD9rwMXSOu959tsRdcmx5+s+bz9QJG0n5rn4kOCD
98A2yyG3PUSOPVwg9+w5vX7zph8GujgCo/k7xL5nbQ364Gkn1FZY3gid0DygzgBB
CcRsyLAAsg2mhknw1/kclDv1LfLEtXzZFlCtxZgjIXZyvPoXcY+hOEXbsmGbr/Jr
TmxrnmbEl9N6aghNE7ZtO/EA1GehX06jn7wKJNFGDP9gVB9s8ZQDPoJV826cKlGY
sW2ADQttLM+wiwqfLXZCmCvkY4MyPl9zjcrAYvCST9vdYPA1Nme9yoeeAoMyxGCP
8PC/ubpH+ful1uCw0A2u9ooTiAN6hS3TNRm0xOCLGknzqDxmfNsZ3xw/ajQpYMrd
7npfFTgjJQ48+Y1s/o88ZjD3S1oKR7svpXfiQIV5O6hCjzPG/qq/XohwfiweavU3
AFUnRP2E6MhBA7jeOdfMXRKDfwE3g6kGaKePU4NTNLMqcOZuEJMQShW+lEhlkKbY
k0ZDlvTaCkgfpyE4EvpwqX6ebsTDyexByIfTsdmY8hlJqq6YD568gTKsR9IryKbm
qtMWfQdoeWx0GpJ0HoWS8v4xPF58d8ZRluH1YGWrx+u4rI06fRltUWW+0IlQ9Ird
kfNV+a2jUjHBwgRExR/mVfzyqAIz9Kb+/MyAoulEp6r4Fw12dCR2BDlU7sQEuEPy
Kq3RVlG0VYcjgzAsr+BGEKBGyTQSkauK/cwaPiEq0BPWs2QO6oIZuenNWl6Tnxti
gBGs+xYtaxoH4Pl4P/sO/WQBJHOkpXN4HNDTNh1ANAInjkAdeUUiUr9eJKiu6oRy
9My+95pdBCEpjHjzfoMyqjY9zJcoy5lN91tiIKXoFBfvt5url+Qnmds6T5BIrDri
WKVBFkcYS3CuTYh26+yXOWH9+IYmr9nNli0W+9tWbm1ZLdhJkzQGEUtcfk2PMNC0
axe6TZ5RjXFJsUvXLGp7q8M0Ll7vSHTS87ouLZsHbi7Vk/YJf4pZKQNPmuyB8O2R
0bTfmaUHpuWhIAJIEo2Go8LDWxoqqfya92kil1DSy1qYWFIx2tNxrQzEKOnuDY0H
QXN0bVlhTM+vQCzvRQD5xyKdI/Q4usHTJjDBhsoa5sfg4TWdh5P2srI/4lhd5C9h
4Z9Bd2epAHX7REjba5L0JifG8nH4z6qghKy7eLfMY/ccbYp/ij4LIlwZi7cUzXFS
OK+6W3S94c1FviOIOK/hH+RP5akCz7ZwSoC6APiad7g2dkgDhTGg4XX3xdW+QbCr
fJj2ZdWGWDmpl7+pbG+50MNv3o7nXA+FlEwzcEEgAH/Xk5aVMZDrglImh7B+Rlda
UaR+LkR0Yghxn3BITUk4SLeZwl4/DOrLcuoYdzvjvor/+kvYw5NtN6iOgvwGsKiH
jx9iKgWUyP+r4/vtcBqkqqenfcAoqVeEMFmx9iENxQn7a+Ueiim2zvCUc9K5+qU+
2g95Mh1kmDaEmQZYNYCPfuQ7iBbjZ87tFhQ7APDNcKeszALWrgiAAH9fhhXeO4x+
aiEJfiiFqojVBfUpUtNBTARH3Q8TmhVmYXJPRYhJLLaEDnLyxVvX69HensAEUeyW
gidjbJydajBY+Fht4yPqp+125HlScgD5P0aDj+ssnhbJ3IgVjuawDuompoiRBMQh
YRxREirH5fWRcc4YBMrY2G+VsW55/TRvuyvNI6/8wQa5hDrZ5r0/5FG0ZfRU/be4
HCxQ07LRTR9xeKbEugE2BfgYo4z9PfCZjjxh+MjpejpOs8+/kYXCGdQArb7XhjGv
UQC94BoL+MkanDUKf+9GUmGGq9+hKLZ7nDqAk92Ne7SvPAWpsc0PZCmjniI5PJCj
IAEprVCTakqLodNKQoZqpDQ6j51A760pJXg2Qq+Ouu5/c+7gq7aeQFqMU49WcqjK
HF7HZ2XjMPKrRfq+KeSHOst/0JZ3J3uoDKVYdHixn70NbHdfhXcqqP9gNGgXvS1u
u+pAgi0gNSzAyu28AxWubhQBMqGy+F6SDsw6sM1fJRXVDfoOl0h927sybt7aW8Z0
dWU/oKzfyrca6k84tlAR65++osKgnZoqC8vKD64Xin7Q0utp1o1hzjBHKhU0qMKh
HHqDoMWSt9rCaFLx8OHtShX1VH2qb1am9MxxLnY7rwMESpO/+uC/sN++O2p0RMpI
WuY+1CQGxGynUeNMEN90N9Bo+siiNih6Bvr2itcrhRaZyjXVfKdRZMVlH5g9/EVq
xXtSBkWrR/HutHjUY+OvEXrfzH3YhNnp6yyAMjTi/5i/6LrHxpmAhLx18DX40hxD
vC3M2S+r1Tl0qqeuxJy0jdkibaEepHfMwZlYL6fpn+ir3F0/N+i0neKZ+xH8jsso
JI8Gr3rQrrn7JTx/opRhBaYBtgWv9SQssNAKzkcTOlhJwFUgXdYV0YBuCvcDoKxC
vPda3kkgkMQ0muvI90lwy3mZXl8A70TmjZo31wKh/nGHg9ljbl/zl8tsip/HWU7Y
Bra1zm8oCdqChx4uYJj3KRKPwyAZ0zCjI1w1S2y6YKtXJtUnJ1aO1IhLdtJdsvVi
4rXVkhk1FIzLg+tnxauZMzkCVhZEbEw8Z3W1jfn06gW+LBf+UpnJKgkD7v2XniEQ
HPEkUpJzPP7SYVCAG9sLUT0WTxaD9WgoOYv16OwRDRZBpTxijU/gH0VwFXBCcFSP
MNUM5vHOsOpdDiopyB0m+IrPfcxZDa66sh4oNFZuMpE9FUwDquQSVfjp/1osqymF
YSR/oEmfaqCfvZisf3S2p9zoqckxusDOggIsyqLVb8SEKlT3ItbQv2H7zbFQFtOE
2VJ5T4kiup5feqjMkLhaDLC/JuFZhFGDAAb1Gl7yxSWGiVWbl8rs9OflA343lk47
MmDfGa4QAsH0kD35iYgJ0kUVRuTpWaC+iaquEL5xa8qLXOF36YeHAZKwlcJTZ85F
8MeLxsCOw3XbweFD0JMbHM5LRSb/x7HM0UIK30qdNtZobKQdzp6q8kGpzMx8DR7B
ZEOxy+0CAJPQuXW5PK2flEY7lLJKOhp//qvF+z+vtm7dMZYZPZbMfKYSJIGWCAwD
1FcWmYMWoxBLkGlryFZ6oSROCt6m0NgVmfPB3276iP6ZNHW5YrPNhNeLpWahRkg6
ZHbP3NxlyLvig/awsSSdAXTdCIJ6Ck/QUvLcefQfKUiWheMnOj7pQnPtpk6MdQRy
9/Xodxu4gwEEPDg5x25kl6w+0p9ttYKmMBtsrN3Qr/bcB1ZUuTOe3z18BCRy2L7H
6fQJgxW+AE5xSPT4+uxRLApclyZKFSSgW66RH4OhQ/0MeQnBHCz2MMtEIrnxAms0
5WGrnGccnOgfGy9BhVBHeYNbi3FVvmDJVNStRvrpzIqWbocCc/iAaFrdz2WUcFDD
agDFrm1amkjJf4T5ddCeSzyhm+dck5lPWiUMSrzSJdNv3hzl308wwYdbufDakL71
orpau4hGzP6FGIY83W07sQ285Z6HMOwRpLC92TUZ76dthFYPURMjaqz5E9tET4dH
U0tp97qmfSeTvDT35LchLIkpzOMhYpgqh5D1EcbItz08zNNObg0nvgjZfsa8WM1e
70IvuaTev0kvaylLvlXfVL7XOYYiAxAGQN4QE1T0yLdyA+YwS8iqmL7RFwVDuqf2
MUEJJPRUV7vFXJT+/RJlWOjL3qk4BZLTjv5zlPgJr+JsfgnqUCp22dliB+zToCsz
KevY4ehs5+9N2nD0ANv76k/AhLS1R+RqxYSzewZo+p+RehHvECvmWCUTF66f4/Sb
4zS025zfr/KjCR9q3wqIMBeHIyFjkAYjaRIBwLURopFWbSqT1PXtZbdjMssQbMPP
+bR4YTRgOGL3rMX16grc8oXfDROkfyGToRuQ7x7qRikraW1ac9Zg+fuPiDq4W6aa
bzj4PtV8l35zlISJl46vJBWVXmiOsDbfIgm005oh5DihgUs8M5QXh/AnPKvaMk1t
PYd78Bmrz6xC/bqerGeOLtyx539UtXv6X46/PF2FqKW+1dPJPA7fb6AWYdosy94p
qsLAI8ENAeAB1RsA35FNyU9QVfcPJQxmqiGAZiXzBB2qnoQk+EqjgWPIGpvTiJv/
mot0jdz7Oo9a4/Cdyfh0cr5iwPzQGGRAuC3BuYE5ay1xGpia8k/Xvdfv22TVW8sD
BYTh+aUKnpqAQkhnOiwFZFHTS4/ppeeZjUbGNDuTJ1HqzYqptZAxpgRb2Mi1/QqD
bCfSp15X0LkoeCNFwWTi4vxZre0hELxU/tKXqJ/psxNKK5TIhANk0Gp/XOa1mqhC
IWgAN5BCRlYyVQCWc5CPrTnsTuWX4TTPRyt7RJkA/HMUrChz/LF9YSYGVoRC+jPn
ZHrjDBfQx7IaLUDx58cR+dZsuETituM075b1MDE7U0bCkZDpzUjGOBG1BZox7vNm
sVReqcdGSfRbSu02RvaSxOyyjwH1oOHi/T4hSwJjhSrzQAaQA7LfykuLkcOQHBHo
jFIX8l7BSQqBaMkGBpfWMtY/glCQluvucXGrF/VbmKTXK7dh+qzW9AIof1pGqAiD
FrkHTpY7jW0BFMszh1RPBJ7tAcxBvF+jqHBPWIQWPB1akePJQ3uDUFLExrzItIRa
p7ySz91e6DufwmS+TtZ01Qq6BgBnq3gwkbZ8ZinzkZ4xexCY0gHFV6vSG3NX5S7m
uSB1prwlEHseJbOChE4/4NEMdJgR5n6V+NhUWFsdUX4BejuWz1iERN7cWdLaQqTd
/Ru3EqX+o94u5jfmtFguag617gypqoKCCQFwLZPknVMTsjGa51+MGF++wWg1x02G
/dzAMVvBklJ1uoIoaJ+jKcw9ccJoWkwf0Dj3pA3kWk3dSAcg8d/HAVITbJpo2hZz
T0e7QVSYqJZ7lQOPIVukRiaROcJ+CrDfSxM3oAvJhsUfWnCKqEenRfOI0kq3CjWD
NPsrbqK+6tIb153W0AYoU9rHU9s2x1U46nh+SpXebXTwZWPCW88PYZMq2QEBW+WA
Azy6y9CxSkgD2emjXQbf80hA3bpLvYYsNHeCR5pB05MkdKZPKmnaS2guwDxwRXEd
TG5L5oTpNIBXm99DyY4JCK+ABtRwQNeG5bFKzYIcTJssizITLBIzfYcxN0ajRa0M
hDKGDV7jBKFIi8TAlZ8eDJYZNp3MqJ5pKtdqr+D79tGEkS7bpssryfIxMvvZi3sG
yoPVp0AqgGHvDP2PosG2JGjxWyc7mT24tvlrDIG9KaRjfTMUKrRXk4rZUxcO2LBH
bJMtecyaB68rshKyCP8yUs3aYFy2ffRrv1tTE87c/LkdRASnhZzP01bNlmCjja2k
MNdJ+L/0ToC3vnKzZvwOZ1nv+z0pYp5KCt200HJuQw5tSH3Jrl45GSLi+F99ZTIK
RS9iFICyfH5uEjmuR5KTpWRRAuM97JTFR7axhTTgYToamJoxaXqpNVfkGBW3A528
PkMrLe/uQGSZPYGgQAZ6GC22jV615T74AwgfXcU9Q6aDaN4h06qlpL/4QxckD84H
hCCwq8iq1iG7yFMJnBm8RIqqndOZMQgNKqwaYEqVh4BNTEut09pJcFcy6ijV21+M
tXcqY2ftmSUzpZNOki/NajRG7r4uLMEBMOQGX9eoWImmRFHO2uu4/6xSKNPzgWGT
5bPyCKFlm73Z01F5PeYaQvOm74xDOA7+TgHb6ZjcQmM8gCMxH3JTcoiRdxXdelzd
hLCyEvlIv+rypv7x7bsVo+WFdSIWV9Jq5opK+x/28aR75bNRrEzQW+1NhntdNPKF
2spd3OlB/L1Yi280nmRh+lK2qi9j7WV6dk6NOE+o7D/Li5KAdRWY9LAaXp5y+pZA
kSPU/RZ41iaR0EZYlwQvnlEuCkKs2KA2dX4UagV/Acj1hw3SOlQqDz3bqHsczYHq
jNCz0ER1UGnk9Y1Ulca//qCmxSheFOJgtDREEEKMLiylvv0XDQ6TYYqCh6slZ5r1
8I7o0qvaIX0R38zbhHAfV6fWECb9RkC4K8sKQndVibkUXe0MQ/R4QozATHpLYTO7
xK2ywIbNb0cfgcB39UdY02Otaq93Ag7ThZKbmEE5MNqtXSJs65oJha+mwiT5PRTR
d9fhAeodlHgCdV7gvxCeTiD6ZOi+rN29pyTGXlbS6jXemXXgeW65wejTD5H8wOm7
hbx/6E5+CxGXa5YOdNffes1cMK3CnxXZnKU9N8euL38JNetI/pphfQmuLu+hr/kD
r5gfcinmJMVwSPVMlNhtynCnPRt7fuLQR9s2J//xhuLVP6zMOAsSpPfxJaIbCEft
l6xrfq3mrWh1H3asmyxeTy14Rpv7VYYxoBxeAuoCfRJi91klujerynsdsvUPCNRW
ViA1ek+ZDHp4CHOmqj/L1VmoXTWP+/ENA+JCf61jfrlTYT99kYml/BgACDwz7d+x
REn9FXRAj8rMDkT/nZlGDE57GCH5+oBkFn762oGmGB7aVqoUCu4A1zjurV08Cnci
ji7PtrlPgmuQLvHYJtJ9+JmdYWnK+rq+oF3aUmP7C5tDEubig814uwFUnJWT65jD
5Wqh3fTebREADDD+pNFxVbRwwBctkNTyj2cAvyskWPJU5tJiiMpmOZfCeXYsGsLk
eZCwd6hgcHfJqCqN+lbaJaOU8drXvWBKetrqZRLeOiKOupaBkybh34nIdXHYU76H
9mFyXAT4KPi1alENwiowM8WYuamjKpAN8qzTqOn/i11ZR4foHj4reWawpRBYnPEx
yyaCLQrIDrilmgluGGDavixGwhjHIP7BmeWNZMmT9euA0/DiBXYxLGJkhBkqZlRn
NyhgjStF45eVHv0SQzrhxItoSiVaCUwC9ko/qdVElQ3DMTcKQGGl5P+C23vwSSBS
4QIOehCtoprOfTkzTcMHmdye39afWPI1LQYIH4s66kbB+ditXT7XXDAyonyRMIeL
PGsQTGP+8Qs6g2khT0TsxDSSYh8BhzlM6nR3aduI15MmkR7H8rbz2r9ETqvOAZz9
9mMbAO16/XEuak43ajsOKmHD/tJOwsD4DYXKvjKFF5RGkParTAePSGJ/tMkREFTI
M+C/csi6ENjDVWTdereRhmZOeEF7J+Fb+DsoKdnv3QDGT7nSPPvObSG2HwmrjtIa
DDnAQhaCvoGWDPJ3Vh4I11VYmgXB2XBTDZk/wxKTwoqm3WgG6LZyOxL0SN5J4FFH
cyhJ+cTI2OojKBStnC0Lua2k+bnUydWeapJfYKRko8WfFYMsZ0Oqk+io4OJ7mC2o
plUcWXEVN8G4S+CAn5Mvhw0Ckyzbx3CILIGePqRm4wukY3CnFLRofY0hnufsA0pB
Q6oCYadwcuReeAS1NiWWGoRF8eKj0IRDOvJMOmURD8V9tLqXWEsux8znDXovYGmB
IizQOo5RDeW9NQ1wXluzk+Wa9gNG4Ra4FZXu75nSq3ZJgzjOZJraNPi7loosqZ/k
nklbkFbwyuURkQr4vdr+11/xHhGS+YZyMrkFujL2VI6T5tFODwAcBwqOZI92mJyu
QakdSoGp4xWjf7Ofa8fS+881+mv16bFS7e8K/VGzYX3AJAVqV3BFpTWudQB+AaWG
icm5HZOwsiUW5bwrKGA6YGkVVDPj15ayAsU7S7l452opZWPTC/h9cuNs/M29wsSn
VXjcQ+HfrMLW6vopMxAmAxtw737iym0lH8WqCJi4WUo8Wj1O3xxTNmCOH3eSwcQd
lVhhKbe77inDrQTahVRTf4UeX5zjtqh2bxfvw3IVRu208/bJLjKAgxROCStRr5rA
XDiuFN0pEFnoKioRjpPV9FNazQokP7j8BlMA8UIDvXOTY5WWaov0vj4MSWsL+gJ+
U3ed7fGwpDva+FChxGggHXRXrxso6isqDNdZhmKXkDfk9QUwrzxidN/SPWw/dRJQ
umujAgM+4spZp57MUgJ8Pbif+u7Hbd3a2R14GsVnyq+LwwPiMJ5fd/5cp42qfXT8
fWMF6gsNMaXGR3sNrxI/7AYrKqsQrFrLDfiODccTLBy53op8PBG5BpjfXdJDfvMv
4O8AVemlNxEOCIvbEbLOUn+AwuIK+RNpG1dpOqhZhOx+l1I7u6vFYIScae0awxBD
l1IW8NsxNHDeukxyNsBSl/twLQz+xLD+IwKgjDUWwZixU0wmku4rZWf9paXxU6i4
qMYLH+wz/EnW3+RwmynTFQjUc1G8EOm0NUN2f/Ug9pwyUWMTG2tSh1kBgW9MDuE0
kGiJMtYlQwBO1zC5v5zZOnQonhpkOclbq82yCApc+tTE7jlxzVa4PuZSiv5SZ+tp
sIlo4o06xjLzjKF/dZAbLjPYycwYeQIgkOX2En00M7kcsbF4Ss3alfogl0vSxuW7
zZlTiCHDZlZjHx7ZR8IefFxw4FS2S34DbhC00Hc6xB1pXWUudqx5kDHtuIjPsvxY
Y5fZFd2q9OQlGdkUNI6wpm11Y3XwBQt5F68Sh381VKXx0M4lEoBakwjsg5ADAiHX
UYV58BFDm0dW9caIjzQJes5OclEQmkQFdV4RXUiZriiVF9MM8cjopwJ4wttSaGx2
pVKLXjIPsG3BNeCTsGyoqD3XwXQydVY/0BiY5EV9HXzLWj99pqb/Q0LM2dAA13o6
IMLiSh83KjxHJBKSFug5l1d8tm9LlGQUlE0oa02q+hJJox3v80CrMdt2nmxnWCOZ
p3xQEh9UJEQ0gtjddVxPeIMs7w6YcspaVL3tzy2b1PWo1thQ3Boq7wE8fOkjCN+n
qo6tLRvAz19A+UMWvpSKY/qHAJGVAnXCB4eEH4kEnIH4XBotdgNlB7LKSa+o7AQY
nuC56zuXxZKeXeojkMZWJHMbhB7ZSu2arp/7kfW47XzTPgo1N88xhNzsvAW8WpQn
J5t2OYhUcPDomN05rJzByzX/wGalkb4SBNXnZ0+73m3Hgs5s18qHByA9B1NuiJ/E
hkl7vdlEb7exfl/q+ENQMlvOKs524ZvNZhdxBZ72k6AO0SMLL8KATu9TESdzj2fy
8WJu7p70m8qM5LW2AqTGCsXj+cGTk1I/TDhMNRGrhSRtsYIaeoYg++k4h5Xez+mD
TVZQZb1g+rv1BU9FXoqBBFEeKdH0n6v1lZnxoepmBgHQcRmnT65qLhr5atxTZw+Q
XpozjxVOOD+5BUWOXutwt0LMNW5yWtNyt8YVHhDD+Hd/CyY7bpJRaymj8gQp/0Nv
6LdZ32NO0OCcE47o/8sR1msxJ8NRImVAVn8I6p2fIFERZUfNUfSn4kszUVMtJiTy
/4QdBdAwbXifHhd6v4iItRLv6VFFvsfjDPebbxsyoQ2ucW8FQ4YiKOBw/djTXn4q
Cm9qx2qCwWHhVI2CYhUSY74vHtRsGHj+LfHTBFqlv6BgHJijLfVcTFtljFPIqst9
bXafS4GX0vQNZm8zFJIHMmD5sJc+M6+7xJiz+37IrDpIRz1GXjyX8gM1Yj7bCAWM
qWS95mBXK2QJ80M68CEwmZVgoWiPpjzRmzDzX3qG6oWpl9/7I3gxe3y+waFOGihJ
7ceSqd7ccvcdEEQH0iprxe+miPThD03YW5BgA+5fK4Had2aASwufNDkGHHdl9tbg
veqY2NMcfRqVDE4aE+u/3H3n75kKqYmttcmZh9rSxo7kjE9gOdxPv9VBMSyJkYzG
a5B6kw3ebY3qk9UBnr4lc5+AII+6OTGAZAYIH67IRCsKZMyJUAw3v2Sb7fagI8/R
ggoeP8Qm5Qya8OpiAHtc8R+cR1lZp4tSCu62I+zy5gyTp8Uo8nqnQmqnMz/mtTiP
9lwVSJf/KDR9UItoR6eVF/fcEBLJRl3JUhKGJ/IgrMcbAODIXoOS7XCLaNZY4CeT
4fFHvhXnfH+HEbmW+l8hcNy8d/4v2UzYbmcGuiXohdJLzXVr4My9Ll81lQQ3N8cG
lpTBb6cMseAGbziUvnkOUPY9bbTjQqT8+ulYCXMjOnFy+bqhfDQUu3+qZ5i6qp2F
1NVGUfH+Hf5qimg+4V4hHxISk3+oq4qohUn62JqYEWP5CT9uwlbUAYnovdPsNtlE
Soe6AKGp1db5CAsovaXA0HcDA+yJz5RlQySji+oq1t7JURLmVmUhB25x6pEATIZ3
kny2LLofmwKRl5U+LPxNXTfSGaRMuvP8dsme8GBhCfIr6T9h5SKjug5BigkFX+Rf
sI8cQpYRimsPRDC3H4AxARcpECVVCG5kLAYBzNLL6CIbajrk3JSPP+rKxfc89Dap
/PMqxnEUJLz+w9gnOuQ5FCIIYiRH7gAHlRQ8lBjUbZehv1Xum7DRs9+7ZlasVRSi
JBx1ZEDsqnh/vHWKO3EpIql6eVXLmlEy1LcPMFuRUzCnjHGLysPdGpwIYDcHOTLS
bOtaIrXc2YUW2cEx+HT3vcb/J4Yi98oGPSEwGGt6s5LI+SkpJxu3uJRy5idjW3wW
HYrzvJQgFDpxq7eOOGIIxWV8DTC05kFTF17kMuHomUK8RctPfCsxVDrp8hnMmhI4
ssOHyYraSBnVNKM39Y2e12BQOgC2fGWS+dPHbR5Q7TP42RcBJUBDdYqKz+OQEGLt
Vo3h1FagO59xspYCntUf3dFgs0qCt/47Ywc+G236z7x/KL/nnGVh7wtrie/7ZRGE
uVAQas3hYKjXsE+eO9Zwp7pr+srMiqw8invlcwjdJahEM6TZtvt/5xgJ/JEg3lDQ
SON1/s8OhjTY5RktgFuYRVNRWWtQGQhY3Gf2Hd+YzQqk8qSIGWcVZgH0hhLXDxQ5
/9pM2GCQPcO30jJWDHj9sUlDU6bUj3YV6mCjcQO+5bcpOv9HnLYKZd14/toF7PCj
7azXfigPcOE0hvgetg53M3cvRm1LsjQGQQsy5c9cx1UNcdqu+muSMgHkLMvON+5V
RWV9dqC8Ls1Y5v5z9NvEX412NAppwayvIKd8MBHLqOahwTysPOxaVpTrrPQaFtPp
tVWvlsCZ2ngT001aQOcMBAi/ZPBG45BKsCWBVE1DpuG5JeWaELddmEdN91pqIpHp
mwpHUL8OuZgg7x2GWeSYqM8EyJIs9ZGDepBm2jjW0tEflaQyn+mA2Gxu6qfMPRhQ
CSPoUtwsKm8ZPIrpafm58NJjo7c3qH2T3uRRE6KyMYWcj442fjqFR7I866sZu2Bn
C20I7ZwDcNhx7RkO1OFqO/KIiGWyJmLzHYo6HgrTr/mDN2BSbK15nlW7B36V9lcc
sJ+AZmbRgTM75xZhEfpVuONhtwqCDCX6IkjTVN4Es52yVnLrKySdmVuNCtqT1ayh
o47wjyFVrhzZbUwwfMrynhGbAjqLinhLAy95HcMhTCt/HpmmQOH+NezJGpGVpFH2
hAurv+FLYWsAYTmVgU8d4kx6eq+CojKvxWd2ElhVVc7mGeSWBXgfMmkwuLFr6Z/M
BHCAv1paBLtnr9w/HGZueYqgmPcFFiiY/K19Q962cn8W/YCRLp0gJQetwiqi5M3l
eGDPX9/yspj77x20i6IVqDL178KJm3yF++Ff7J8IQ3MtaTFg6HW7Cp6MLYTzme2C
kRnfZ3p4uWP5x1d9d8fNdF0Esn/AdXQWA2HOU7e6ikvDlXm4YuzjZx1L8U+UuKIH
i7Doht+Jf24eg0nL6UfzPwRjSdqQduyIMNvbX1YRioQhj9Y60LboPN7hE/58XMFm
ukTfess1Yxk0QUwig9yV0jX7MODvXYqPc8MEl4XCHLwk2s4882K/SvkNqBePKW9B
AXVCt96tGwmEfCS9xuYWUAcqo13hpWMgrFoqxwJF2WhBIXtuW/gRjcCQqSVd6ykd
UreZsHE4jDMNmKENzgl2T1a5h23cH+bIXddCDdfAdtJqz1lu1eZoSyUjkmL33NG4
Nqkl9s1qyMTt2W3aaJau1IkNzDeU0BbyxXaMTHPwd/NfqCTr3ccvxhwLs8riip94
QTij4e/zSLtM9E3RctoBytZ4LAK3RNVXomn4gER54u/HFz2k4KVYxW8qwOjN9lhB
/rZxuL2D16+0Aw/AreRb4D/Az5hDza+b1sPdyMEJsRq9wFN6sPbs3hU21DIt4Ub5
Ivt8v+dUvDQsIQTLOuRGLOGcz9DOdYYUHSFY23Ik9rxZ1lnSMVnxJ3hbtxxL+VMc
6gqS+VuRc6aq7UwNYB9g8C7W1/jf7rgzdhGxjwM3e2LupQ+D/dOTBfQ2BIPJePMl
h28zETu9TPMJ31yX2xHvWDXK2pYwBRCCn87HNKT7DdCyBv95jOlCV2ahACGJmRjo
1FJAv+tkr7fAVGpcibG6HqoaiG50KaCI0upToL/5N+1R19GYujUcvUajJ0a5si8D
6Pvs1KXjZcuSAcjIa5uPQMNHVK87v+jxy7DtvSR2h9NZSp9uTF7T9bObLJzmaLSP
Xhe0aqPo6TG43iH9Mg5ie7TLovTAKWZ0A9cpZN+lqkWMQSoYvWE5wbEQUWDJvSYh
wtb8YPAECXTHMwFxAFUITGNw6dyKPnmhWf8SF++2PcsHAKrQOEpRsh3wRhtTkoYJ
lc7/KZ3Pt0FuD8D6BxL2AnJWuaynmC6HK4re+KU/NxeGXJE2s25VO+lqYmBl04Z3
hCtExrXv3E0j7Iz9wHgzuf3VQPpdmuhro8lpY1fDClOP2jefYrORyrdnDijTHUc/
kVd793llNNk74ios6hXgr67ePTGLBbtwBVzJqcuePA8ErTtAfAp/pSbthlYHpNNj
xWN3yy7bHRFNQvVUR+8MSNk7uVvbhMs6fe0VVXavyAEnMntkeRYTPm3ZvClS+LI4
wZzs6pU1b7D2tnZ3a81UekUgpgBwkkxgIxRvTVAwjwRTaERProBMggimeP0SVHtv
HKKz7f2vDDguWxiczzUc0Ud0i68l3Z+aTYa04VIv6yYQ1yY+HIz6STzbBt+1BuC4
LpEtzxDY+vonye2+JP/GO2pmImqn0y0kRBQ0pYuXiBfb0b0iIauqimFywD6EPGjD
Uo7E98fdltWSrdnnnTuCeDuUHm9bx7iC7+egK69RZVeMo3zjda0nWGQm2GbQtAd8
rnp0PXLQgk9z+Gm6aAHQy8WTrpIMEg2KC6L/y4a1vhwT9FPktZOf66L0I5otn6hl
cBoFJcKEtjd7aRDB2vTgXX6eGTuNeMlKms40d63fX3rPVjeuD5z0CzdOnAitYSjZ
fXrB5sczVW6XAt0Qs8wM6lHZ27QOZ71yIYchSCvv63pT4TaObtoTrVbL2OChxx0R
3Sb130CYOJbXc6WS9MtkCDX1skgw4Ke+S3bZGN895DZgjLcSzp7udNaD8cu9X29D
BHphbLiujtRRjkrwQfGjLriZkwoqfSeuoduRujiF2oYr6B4j4xj2lUaaUVSfY2pr
62ak6fhDsUD4nDNQQiDh6MoaqtkoizO8sDNHDM5aoLG82WK7GCosyJg1xirOoBX7
WUc8BT0RuSxxcrh+doYYn3Q9+ArqucjrxOw9Ib3m2SqThdXg6/XV/AuS1G6eywcz
8+SNv0V3myzyZUmb7NRyNlEgHYKTfWz2tdYAk6z3ob1f+1sr8CIy0rOK/+z9Dkl0
ibhI1onAqbO6m3thk+Ec6bOAtjdPUt++ntCF7gxRxeCNO32DGHIXXYOx+lR+6yD8
KaV/Z64HAGKgTFptQ75LbI9+ZgVufgmckRHy/yAaZR+2cBNQUY3A37r09VKgVO6B
B8Ofww4OGilqQ2iemI0sLlrLA1o66fho5NhcMgfuvFsBp4HeROpLiCgQEnba+Ixo
0DjLvVcLpHnBZcM0jqXhpxiSaczfeRooU1Af/aEuUSNvJVp4imaF4ALsp8TRd/2/
8bF6QDMhUhepd7pYAxmLJw3fFuwXIWSsOJdDVot/lCFSOCChZJ0/OFF1DZcLBze/
VkC/cLvqn7cs51P9xY82i1gXajufklg99K0af178BwYJOVgPQ9FgBgcbSvLKi94Y
jytSu6YHYnnQpUMRI0xtOLzW61cS099Ea9ivcWx7CrhzlSMsxHjDHccomjlov36y
1yZh3fshZ4l6KcOLEKji9C0+USnyf5AgtUHjZ20cTKqb8tHMmx4h3FZm1QwshhNN
Zcx9uLbG2MX++8vK+CL+OinQsQJJADn1yIoYq+OgvL9pzsiNhYpzhrxupyET+yCe
3FNgHwgrSUhVT1cSn8brFebDrZn/hOxgrlDbzRB7L2FzcQd2dPTuJERwatBjeJoH
DDLM22WmrNCSdBSMqzdA8O9CrMqb+xViQJYDWTZqDApVtsygVmkV/fQdAtiVnh4c
Oe4wWvia5lckOk//WEBa3Pc3JMDi/34qf+qsImhd6TQmPcQiG7mB/lq+OAulvZ5m
80C1Z27yZO2siby5/MsMTvMdwGqaPGuYg0bHrzvrstp6NQWG/Q/aix3gSnkEFNsN
1vogtxNDD5WKNCxws6LmbgZi9BhePgT8GQRuzV9U7EKf9WnZXk/wYGMQ1v/PTZl6
0sc1jOPD25147am+i5TgUyhU4w1nKpTYTEHiZWvVHKOtGENFa2Hpy6io9B8xcabj
ByMlVYZ7WAx2UkawCvGJJNm+diXsI/b3g10RgcxCVB09Dek6u8+iLl5TkfdnhjvO
xxP0kjy1NID+G1mjWiaMeLn9E+MqPLbQIoYKoS8ffH4e6bjD3WID4rvXb95dHLbd
I48IKRLZMn4Q41pLIUiHAVegAAVxmy6DbaNe37J6pxL8mrrJoFE9NWR8Yios+qSS
rgG4FUW/TzQ2u0wUB3mNl1uCT0zA4as2kK1JHP279spjbpUl34m78NXpMSFoNCWz
Hz36G19anljiYxV57TumbRkV/1w///4EQ4BZ9qnhApurbnjWBcbIdetECQKr9hlb
UihLxNbe6sO3sl+YD3/InszEB+DW8q/fr/35LDlJzRV3zvQ5J6a/9IO0XP8C0WPA
BuKo/T66HnJ1/DPzpyxngBhmDBEs8U/OPZFhVcvJZVW+pxbQNkmzgrHBqXktqbyb
5nz0DSIiDOQGDI7HdVuWx8bBEyrEJbEp+P1oCmc0zqjF1FrU95HcarBBzL2tY9CP
XTey9aJjM1mCg6lNyGsq6PNcT8NLjNqkQ5C/4pjQnPx9MCgpc8Tk27+7UJ9NyFVO
guVuHp7Tkdxy5EAYOiynJVk1dZi5+/+ZylJtq+Go+BD/tmUPlKQjWJTK2c1Hb2Hc
A97ofB098GyUAIjvFKBYTZaLYLEWdmxV/NkT96uKBezzMZZNnMWakwayVGCfnXlz
D3K/8rd0pVtXUPSgwMBwOAMtRB6fAqfPz/RKtIh91WCSwpwpxvzeXSfK+FBLZQsc
AAB+YtV2KkX2035pRpzzHBCOXOQ/8Elo0y1CNKaQHVS0FpkPK0rh19cFIARD+naJ
N7fm/sCXvT9hxdT3iZlG9kg/ppgmOwAUinMlFIpIpsju1YziM0/mCA2C9e5x5rma
mYg9/hY85TipEhoXoxQbb69xt8glc+maBXQ8IDizU2WFJNRsTDE7rJhhIM2qol2w
8iGenzK3iKt0eIb56c4NTIXRt7ziwVkI2ov/T3dtlEW+NIGVahNj81kcO1dNZhFu
q7288mehGw2+tbrJzwOlVzwsGeZpiDTk8NX2jPYMAE5TvHEEyVZd/tWbN8qPqu/z
QaUZ+PSMFQdkSRmYtWNciwCHBNdIJPkoFhV40RVrMwD9fML9Y2ebB9iveKtHyqji
Vfck7a/KZOXcWSZIIhu4rgXsojp5iHdo3ePT+NLSCcwNmwKifjWuH1CDr+8AlLDs
+rZowpo25+yA1So/WUy5jzTxhoxJDo2fPzzgQmljtyLqGX/pCItEKIguUnFm0HAT
PZh1HQCTYyzp1UyiJiEBuqcukjgUukDVqLvZEu9MzDfg0Fs7LJQFggWWD+/K5+M5
4MaIW6vP5kLP9w6sm6E8CQwNa4KdlgsX37V8ZyZmZ99vl6KN/F57XYQWdgzWuVsY
2dHE5734CAuiGqAHhgTguih7afIAvXpOvmnjNsQ7ODehfuydulxTRUsb2ACuQ4us
4yITd37TyBPB6y5n58X/VNo6z3UVwbdubDkTuzmKwEjWsUQxmMVuDKGfHEe5uAVK
hvclJvDQJjVgDNO1yUhI/0NBO0JdwGA61k1GLiCKz12h4YNsY5C4jWVS12XPNMXB
A+YnNYvDcOKVNqPIiAvawOh8YVMMKoLDdKD6lk2IfweOLNNwjZK1VugadPGZctLt
tvTVmq10liNq+qUgiNJVHY+eF4kR1Byed+2JlhKmyQzkuXdPJBwx8bQSvc9BUf+T
VJPiXgxMRbQWtVslsxUoxd654UTs8nhpThN0ytUisb/cZu6MkddN2iXhPgKBN1qa
dxUEqpbtm2/8YJ4cSTAgUk1wRfpN3p0Yxjv/l+Ag+0tUVMl70mJN4U4VQn3b6yw3
hFj2uip9B89Keivpr/d51TYADYfdrCMHYC2U/HiMBvd9EGQlUnB+xiAYhBMZL1PH
cpxuCJJqN4er0mZqP3z6wuIEcWUbzYAlKymSCfUqfU8NQSZPA9t9gi+hzun6FKwQ
aPK5Tw3ceicfhjCAihV9QKZNNDaG76w9aLTJzwIv3TER9plWpUPEZNtdyxGtCD7T
NIveZwnmV+JHSRzL0cxjcZJq5aLfxzgy4NrlG3L4It33tkbklYjr167e/8UoHmwR
u2DpOMvWx/1oQa1evotWM9LobaVKhTQnQM+j19ILxj9OeNK7h4UdNrnNJIhCh7KR
cHzCk2oElu3QTpaQLzn5N6vb+nlKciEOkHyzGdyOC66uitThXh9zDHUgCZCZP7/b
y2SzE1oimB/N+6zNrNPjG3DNv6UfVOJpjNc2nYHmwSNHJ9gO6RUX76XLy3IUebv6
TvRUQUC8UiQMfH85ow50KkL1tO90NFNdzDYoPLvPki9f862drIBLuweNKNN64LjX
puY/bWAkX+sNra+3oxQ5B8JHJ8Ma2FmRkUSMkwUZdC2XufI5SJHymWeMAa1TCAWf
RzI5RY8pe1WeGpYrFoCe7maKTzXjy5y6a7n4w/Nf4orE8qJprTHFP6cOAZRy3WEW
oxs5MsLtcFuKhPz8GGWnsPyN/FwHr0znJZQcs3pK8NMWEh+cEwdLLh1cHTj+vS5g
tXeihWPHD/bnZBj2w1DY2knLYE7tGE27INBqHfWNoolJ7Mtkivx0pf7Z7xjFykdX
V8T//y9EN5Nj7M2GnItxjded/CCPKLxAW41hntvXgA4Me+tSX00Qr5UF0qUKLyzL
1HylGuwyEF9fCjQJsnquoJKC5879aPey/YqkwN3uORFHvYxooHXWq/Og9Wda84L0
t+gumyULi+oZho4NIimncLxywFgGYJgJGuOq969cLpwk3tuucCftB81+shkCbBjY
77IHvnNXKSdDY5pTzXB3mddNYh1OZw14IveH3p75ZjU9WQQ+H8lFXPjovwC2OxNj
IgMEiOX/j4hhKrb89E/IWKiadjyUHfeC3xk+LfFKqKyaPz0VmnI+nF8LHkuS3Pcn
3u0hluwFQZDAYvjWVEWNK+CQVyH+Vs3o4c9EDupku9PdDpIihH+KepLmUwlzdzHf
L1kFd/D6mY/4m8cs/NKUJLSfzBtXg5KmJYX4wYR6ATVGNa2sQDNrLYBVNQflMiU9
P36iHdzmaJ6gkl0Xo3wKVIcLM1bXjPBO89UjkEP3d5w4w3rYNwrA1geWpUBJ87K3
e2bxBfrxU25hvuMZocO4O3Yw6b2FJBjwqIl7dY6C0Xd9QvfWC0/YcKAssmwYNzqF
V3ffGsOL0tmcHN8p5peMP+5DX4dFTiE+aAT9vifh42Zm8gJQMnWOIseedL4sq1g3
y9KpB70HgRq2tpVRjXI6g6CZX5toVb60fvQtnkHeSBTO9SMC8G9f5hHHEj68F18h
55x+V962xaOyJJdTYjR0MhnDkMJI4GUW988R2t/HjeSD0OnfzzD/VhalQt/SGBtC
8EEh+s4tPnyVk/k/6XVyk35KPllGjCaBHGtnCndpXKtqJFXpsa3up6GwNBntlfsi
2dpswGhISia8LF+XqrnNiY3o6NyLumJf4SD7qnW53jHvp1r24Hm+7RpXn/PxPW0d
gU4poedHEZu8IydOZanVb3R6wUbK3H8vhAvaDzjeIzbfBBapwyPCB0B5QeBeqLfN
nPD+h5QNMOMMLT2oYWcpx7OTKi0f/OShUVUnV6iq5/ud951HPlT4MfO6B73y3Ofq
uLLnRRJ0rPTkfdK3+xGxQXImQzfwwA5WnDMg2UXf0gxGns/+fP3JzdAns3vUYiea
3jQQWwnGFRK6MPKMheenBC92jq/l7gVdjCP6UR6nd/btuXjQT1ZgdBm69k4JASVZ
U+FsGDYn1pSaN5Bxl0oiADzuVkPsBe+bBXDuJtCCdwqDSUJ3OYylSDSsmtlp2D0U
dhWrF7RK5BI6zrIe2T5+IBqnZapc7ofFIm8+wBaPLmY0aclEcFuH4XSjKvOop3mL
FugcNRC51HqxHkuKRwwiqN4C9yX9L0Mo57v53kZ/f0jY39escxRXVth6bPjF/wV7
g8TyMkqccvVbSWALSmiJjSlyF9Gxep2BRk6otn6l53trbpgntyEKKgVtl+lTXczX
iaIz2HkQHoqs2XtxHHacs9UhCldEbvLJtMKby4YIdyRK4/bC5OJ82VHVK0PWEVA/
bUiTA+50lpw7wXjsJ2YVqUUz/woJClfaKw1MJRYsiBSeB/lr5G5x10T7p5H6xVQp
8W84+HTW7pV+0WPGvuUai6/o8f+p/n5VcShW9HRTk4PB3eK/eZHLZftSZKs3mJ5r
63e4Aq4ITsnkWfuU+ppnvyLAw+iiUgtHVaoIOw433MmOXp3WNZd2UXLjrXQZVTHF
yhhkZIEAE4i1ARcRWqdWEgNHZuRbs31PTPTltJTXypp/G/GAzfSYHrjkz8wYYN61
vsU2Xl/05JNqE6XQvdq6BPxJL8qEONcXtr7e31RW8a/hBHfi2s47CF46JAAlI0N4
hVvXx5NS+Nz6HAC5OdHqWTYxkvEzqJfSAnWCuwcc6gD7Z/xMPl1m2JiELDZmLKOs
WDhQK3hsFNN+K6uwRt+2Y2zBd0/melZRrUMlfj9UVpZ+HX2w/ctGHW54JY69JRFF
MpqpFmvgZOawEjW5wra1WnZJPvdS0LOk0+tJmdp2JfHNOTlj8MgPaYbdcMOLTZFn
KHd1A9fdEiwO3br6BV9SuPq9IA/VDXpL4ssQ0586uMXb6lTOUv9e7EF5xcBgQBdx
nX+eJeUT6pVR5Iz0zi2mwAeQSXmt9WHvGePeqTFpFC2AwNmIBJLNHwXQTZtOT4vP
mQ03G5vCNRliff2e02BGDBI8WEhpNUfJdF3a5MiPE0lqkGVMYbr+flolZxpdOtC6
JJ3lsMUH63ljv43Tu1P/sT13byTNSurnb8gNpIpGciwS9R/1oxAdcnej2T+FxTOF
xPJVg4zJkIihgRVPJ5nFHLa8qqfwYpEFGLum3kaWlVKs1msflr4nKjPKzUuyCYaK
7d3pwVeOq0nDbT+Tp3+lXXdolVF36pgw4rc82BKXsw77iuqZCPNaUXoNmseVjdYY
RxXWxMu4Nmce67D91l6vNQeLIW5aZ1auicfSDNegqfd1+eu0gFotFumvrwxDtBfH
9VBEUBic3xzy96yhB5PzM+SuV5BdHtgXduJmn7oPIfZkw4vXiqkYdRfPl+NUXWmq
U4K6jbwZVpVCa5qpZcNe14nc4FHXJ8iinKohvsF/1AceHEp20ZmqBER/kZ0P1thu
k4g8rCFu2SaRq4hgLA+e9Gono4ALw4svksXMal+JmW4ExlHvr9O3WDh7RetoXpL0
mUgo4jN2QIREeFACz5n6EHSXdmCFjHo2BXnj8Y+y/hTlw9DxKsXaY9HK8RCU6AUL
NPkuaRT2YFnPQD4aUJsSE1vcWnmAlhDc5LeAPK5QGtWdWpMsR2CoqcUiMXo6zOIJ
51y82Hbny19uwXkJf8nc/IHLXQAyNociz/x83xsJvdT4IE4u/8KSESC0B35cz23R
oaADGPKwGNNgH5sabyW59Lwl9E3QmfL0Mbvv80G+FdEeyHhZuDpxdBv5SBhSECHV
lcKsypjLJeqbuS3tvP+a+4bsRKdnF2B8v1zEwojcDjQxusIWFDKLdfELrgzT/VHB
L9A4iXg5r8wxlPe6dFPB5E6dY8UhToJlfTpnSOu9OPEng/rpwQiKVtgx6pKDCOXx
ImzWrKRBKmtv/1YNtCjPmSh5ggnQCQK7g9CBwSED86LKJLS/lC49BIG1VurtzSBk
6PK25t6CoMqTCHSwjNxh7pPtU1HwaNLm7St8Y2SaFXf8XQZfO6GKrUbq0MRe4jpE
FnRlZ4JEEdyM6KWozLURavKMWn/xrsJcuUeglhQ91nYQsQ4UxT9KtTaFhrxGOE9j
EHrOiS54qr1Nb32I8f1drI5FrrlHz0wKe25dNuQDLqxOCZ+V2e+Xh83ZvjlfzrxI
zUvDoL8Le/XOtmbLiwpMrS6sRksl+blLr4HdH18wciFhN3Fzr+8u/TlNRkOkCtT+
GKWggSDvfS8/i6FmYgAsMEqAifvykWbYakDwQce4bB5nBnYpELPCRgULgyAd4cCq
vihb2ovrSY9p7A8DDL73Zrm3RS3mSgfha4z2dzrq28Blb6ZIsD7eB1x0TsfEmFll
qZpok10UVYH37ybrCpy8BSjsOf6fEiV3pKkc0rC4bemwBlTXQ5wUTZayPye6+F9Q
e+z3M9T9apQre+MqaCfKY9aOgQszurXsJdoHHpEFXilscGFmTJRk2M4ZGv6a4IoD
fAG4ccQc2QsPZlL6CWrhhe69S9kUIdiJv2Y+JL3LizMWOlKOQAm1K7cv+vCpFZ7x
38/VLYjPfDU+NRv0gNqmuxPUKgOyNAS8b8n/GZjhvVkHCu29P10c092BS0QzdVDq
VlE+S9b5AMThtI3edtWArBg5poQhxBvvUIm+41SQwx2/QDbigJFmr2btZxfKtAHJ
wo4l2Kp9RvO98iNLv0OVx6Pps3Nf67J5yWJ2ePCNCDUh6966kvUQqfnnZUvREdat
aVvVq2yKu+c1hdrWX2smY7V3JHlgnDxb+XMFc2m6TiN34gnxB3YoiXGuzLOK7ciC
xTsQMpSRF3nR0zDId7pIsHzuVXeTEs2WlPqbBsWszJEFdzzhunE42visCo6Pd1Ad
n50ruatYjSg+cdN9wv7usn1IGQUlz8Ja9jo+uHdobyAd1XiTozz/7iJDgLmM5vec
HvCAcLe4FCjRA91VcHBqbTB0hcnvN7i1LDItHNH1bXcSrJM3pNxy3epoGPj5MbZm
aF34D+2GtoCCLCz0TPoO4qU2onne4cLNHRzJ1TnrNogdPqY3/2Lhex9YqloE+pX2
XSvMQbQUSR4b9wMOkgEH3f++SNz4a+NKhuqGwQydZJtbp+PO4rFQw87q4xlthE9J
sgMRDyhO8Ef8gc/HZZJp8w0kSQBfAcIWwwAJPZxEfjF8JCRarmoP691TZ74WgvNT
p0DVDle4AUC16Wa+S3a0k6qkcDxQr6RFwrYIPbbx7jnN1v0GzXlgslxrnbat6Jcl
M0PoztCNnJKbVTFU4Jm+dset9/17o+NDaHw6UJ8S7v5rcZ/Ut+VtLPSbMZQjutry
LgOr2WhTNTyDTND6Ejj4NsjHkrQuEkUMX8qwQZBxwo4XI2ZDr4qq/Hsrk7ZFK08U
g09G745/kWrK4SS5ZeV7/1eazvtaDYUkzhmFRDgzW0CHltAIwaEJ0E6OEMePmVBL
C6PVM5ycv2W9JAAY9g2YsQ9KpnBhsAfcaKSnL0uVxGY2r3FLa2R53tkHt74rz6OE
cizGcJhGE2fqN0QR5cwU11icXPywkv4PR8ECgSkxqnfvZ0TG3i+pmnJAz7xskrNC
qeVLffV0xi8cUN5cVol846R0tB+jVpcLzxtadfaJpTTl2fAet+Q3+MQBPeKZdjSQ
COVV/k2+9ixhED9HGPJtH2ZhWG85wFHlppE0W+6dDRa7LQoO/r+aVuYGzYVHdfos
xDaWpaG7ACUtVDxMCtNPid2qiW2T+0ITol23DHETJXSpXiWrNz28psDvD1zojs1L
OufP7LG/z703Ws5UlUDjA/3cznan4irmimgPnnT06kvHH66KHN7fIhAz2OfjHheD
UdKCoRik0QSIzrvo39oCMkXUiwNtOrnQIvlF1NaK7ZLW0nt6KhVamajwqdsdoXjs
QjV2ObcSUcJ3kDCSWwHlebpH6wByl0esZ0vZ7XJZwkMgM72Ukqd1TzzrnweNlVMI
/84ubwuNbxtZU7azyvCaeT6Cu1/VHdKTfi4SSgBDyTVT8SBCq79sGkdFYZKwVGYg
QGUl0d1WmZZ6eGpyAPYlfQaWEw2XgdRt0is/yU8lYib9rIlvtyZc64OdXtztecz3
eATRcJhHW8JMn0vI4TLgfrChRHXIJ60GcQ3jx8pDiJTqduJBHy2F5r0DE7g/RxZ0
56ocrQn4pZdNTLa04QaLeyc0J0HNYldVDwTNKTjux/V1akoTkv0nBNiza8oJ54PS
8aVmyxey6mXKm5N3DjnD0QbXR9PEHLPquTuDbvyjgUUOOfWsWkE1zHs4ERmihLvo
IBtjf0NnMGGMjQBXGomzPeKjA7k4yhzcs96OmmtrrmOqNvqEGZbA9eoWnlmqvf3Q
Q4xKDOBUD3w/nnqgaRbSH7YFVxXuZ/tYg9MbgzKk/+7jI8KQFZagc6U8rkJepMSC
nVgOEXObtX8qILHTIq8Y3+I0mTdu3ZeENvDBobKZAWNFP6nHYqaQaqLhDIdFphYA
lKUsyeKc7gAh1UXXNT4jC6+9qSvWKdEmv7ThkAPbzu3gs1KvqnGsqlH1KHUwyR//
GCqkz6w7o1sZRut9ye/FhikavbCG4imO/Hxidtcf/1XNDKXZkLC8Tp/tKo5/zZwY
xjzowfES1y0KZAA0WoPjDvOVtzoe8wlkiYcxCODk551P19ZyLnhWTYmHIinAqa5I
C5r09HES/g5RUB5P9pRWo03ah7h0cyDD9KJG7wLgSIvrQnCvpxo0edNJ2S662Vk0
UU5WlXy2lWtMMqvM8ETF4bjmKqy3ZzJ5ISH8YZYG6keZY4NXpO4yRR1jmcmJ9tpA
lWyrZLfvHJJc/fdsnyzC1CXV5W9xsysf9eUNeyKAPJKc4g/7QG/PNboSJOd5BU23
H9HKMykjhbD78YkazrROYGlSn233D3ynMjr3tjjiS+ly/aL73e7nog7QEgIJbfWI
50QDkh07Uxl32wwz5dbLn2vEjN3wmHUCzwKSez4u8dBc6qWCAI6gNLZbgng3t8AF
o/iuYtAm6eJIk/W/IaTNGnF3Uf0+pyY6rrPaYuy1kWpz5nP4n53faaw3K9tAv0XL
Nmdfp8z4d9cn7jnyM7Kvb4G4rq6ivmp/wHruezYTrmbqcqus3W803WiblQLbDLVH
n+sUqckZ9ApQHTxGvGGlrOeOWyNS4L4i+7NhZsprgo9+JFcPT4IRy5Sv49TpNkxc
gQyMQ0Auy3F3Z33wEa47ignjwkrdpSdiIVOx01huShyWlpJ2DbZNz5nQNoOu8WOA
Igg/Nl35MRJ7nsUACjOx27wWlo9CcRVtZYXdX+eaJpeq/daTlLu8yDtQp/GZd+2A
+cA0VH17Oq+hcae6eJDZfTDKKbjQNvB8pAIB5Gw05qTy9ZrTj+cbIGZcEJR4liMw
BXEhcwMLuMqHLSHWcScsLvhKC0oCqK7XzHXAZ/8rl+oWCNFoOZkYPzr3AtaT+o9V
jbZ2T2gh6eyq7pqVXqgkJ3j8V1ojrLvKPvJF0VGhpjkLu6x/eLaHRxO2AnWOGiTY
IojThEwtreQL6pLBqJoWdVAR8wMJwdg7l+LOejd+sl1UxKoNMnl0jaBqyxb057K9
X3zOOKTaApaX+Xu18+wcO28Me6XU3XHNSnDvmDOxDLVH5KJ18viBFymlybTNPBzv
x4jRs4vjjF4dhVR+lc9Hq1brZs3IsVie327+pj2koAK9GO5pnR6PsgRC9UEdD619
eUvKg7tD5wQdix8LgZUr44tYYwEW3QXIqcSVXXksG6yguy1oTJBm2thjqtRfcGW4
3kf/yx3svAJMCsnltWXDFuYjbno9j+k3b3H9trSftAYrtrVjSu3xOYWjj2cE8FJx
ZlpoiqhNgqTQofYqSlPiHDNPT8J3xx4Okeyob9YH/wdJGiMrucJgVJpkGfCPpcrM
SoLBy0ixnF3X+yjVYAdufyxTdh3tx09kaouDrOngP31YFfatGcoMd1Wiyn/V2U4+
JWr0+IxJuAHSWzliTH23eYlMxJRxjpLkPG8mc5wnoCaFt1DVXh9cVe6DS3IX/b46
Mhf0fv2NmKMQ0/IvC2iNhRlMGTZy1ThgjEzaF2ZtMGZjZtT7AWobWUZmwxw8sCkJ
ojrlOdhFg8iVUMPJs4FyETeZHWp2YXNH92QCR6khSzh/BVUqkW0qaKin7YEHmVTM
rI4YfpO/UjiiXKliMF31KBN88tcWCeo2OaFy/eMEXZh0YtfWtFYmqC20aHWjLTSS
BVwK3igyNlG3sI6vaUIvzoC0CUkSu1RhzQ0syEjBsgHQEO3TIbdFIIDGXOmPKJQK
DzHzQ68ryDxerux/mX670RUr6cP1llKj3eNpxRuvnTc4itSgNmV80MR9pjlENudQ
2xNK/vsM1QoO/MezSjL1smx0J2ObtIti6tlfBtFs09w+cdM9ll6bwGTvr2r+zDGs
glZeNHYEcPe/4uFCgR0iEQZUqmeACKknQy5EgrdrJtd51oDsXtI9SgxhcpzIvrgM
emX1CNsi4P3f/PzLUyaJTadnjHda/mBgxTv8lFeHyIzpPwynsbpSfreX5cWMG9sU
MbrIxYx9Nf3hD4896AmXmwY0n8NMwQvS+8a3xVmnfnAIf1++xHwgIfvvWTGjv/cb
N3zg1yUHDpsXEaXTONJVkbZYw7ZS7D+7XTwcKnzRjYyZRIy4UgNsd88bbn/PI36G
JbLd4mXzE10wk3Sp6AjCGO+hQXR+EG1LwMsPADcs+MXiMzTz8fR5FTylkTh2EePe
AXMqWqXu8Sh+q/MhfL1n2trz6bNcaW+3pCkoHbKt1TmCLHReWfvzT57nFGLD5SCr
Un9+OMWWWvAHZgPQ4+sNkhgOuU3eETQz33olj8YUtAarP3fsTCBrpJ+leabfINt7
1aur8qnzyNlWj28YU6ENHeOPq+NtCk4OG4JI5xtNfcgzjVlWWxxxHpqv+4LGZmgq
zMcX2tZcl7eZ8ttXyeA5FpwI6d4dL0UfBUg9Bh+2+SVgcU0WFmL6ht51YsK+3QrJ
n6DR+EK36pYq5UPTy/aKMgDQZGH+rd8/Lq/iAzurjsHQuildGYptoz0nLoFrsnM4
aSBn3xLPKQGUsHvTi15Vnvmj7S0r48DUV7We1r9OJZJ8sKwsVGaR/va211Laag7H
n3IMJoGFWvDgDkiWJ4oIPoVzKTPAubezwAB2vDRjB701eILAWEzflLfK+Ti/f7GV
nNFUSJWQQFJzSF3rxVK8daKiYKmnJ0gwAs2wrPE279OICSh5G9X56R5vSnzpE0Cg
UwPnETqK0EQjAopNqQlwV1pRyhbv2qh9DHskWFGBnhjtAW/FaKw2nHEhBp1vRZka
dFfoaRmsqyyLHAXi9gGKIFfB/CKzd1E55IXQYbaG2/tnuTwLLOyDg+4bwfD+U9AV
a6juS6En+FIoiBd5SExa+nMJXXe9TvF/HmDz4arzUGsRPYWNjLL8eoe7VIeEVHeT
ylh3PnAVeQJfrVxOp8pKCFYLHsfDpcHoH6WzNh3I1J86RDthqMfxHAVLf7GXURwi
lqWFvMM0tA6exxROsIiL5Ty3FyZaGNzrWO7Oe4dMDdseeU6oV9z1eI1VMLYGH/7c
PQEAPNQ1RSQnVGAOxvGlc4Qd5lys86TlRoWy4P/IkUDYlSSCdrfsDiQCRr0RjUf8
rn1kvKOfzsOmR9U1jGv4DG28AYYG7cVXuvlIudb0t0SfwkNcyZVtk8Y7iHMb558e
KUh+hpr6NDNtVRBSrH9V8jIP/HmUUyuvExXcDLRjh+H2SqQycmrKbm2aFFTvUDc0
unovBvlcvMuCpaOEog4207EILch/NP8SqtMrQT+qHOc1s/+C/hC8finTIv7LZo8O
rwkTm0YP6hXs4LLHL8mxpb0mkhZDgUL/veF4lCGIESsOqZEXSe0bZY6Ut46FiIy0
JP7TO4e4a4+aDmO2rrm1rdSnGPlaftSAHvO1NOyBBpwIQBLmGKnvBh6lDXjR+4mw
q//B/HkxbPVQ3UtRv/+Ygbph7tRruQFc93OiHTeEcTNHo2qsCQVPaunzIzXVyHe9
xkhQnJVrZ21gVgQC1GHD9NSls4y/u6pZewUQc1UmDz/fXOyFyzxfp2e3uxl9983c
Ipb8zN5RzEG81kHvsWmgWV6NrYMAA1Hu35wq4gKgQgKrcXR5IYrNHebAZurejRRo
K3PyChC+5dwe29g5UPQGuA4lhu0g7mdfbU1i8r7yZAxMIbZUVZbRd6IuykltLG+G
Tdk3olK/t6jBlbhvWpTsV779JyLDxeYcLRh/dJWjFCOSDbohhyNm9gZ3bV5yhQlq
/RNW71+IoRhDl1PD3dmZJTOfmhirBW25n0HCkTtSNI++e0JtCzCVq8gwo6NJ7knd
PrjPwfFlrWw9pgEbY1ej8vtRWB6M9Lht1rfYlz3V3A9Or7Jkc88PSY9Fj00//LBE
fcVfRPgYqSDuFNI5FrWsGN+LB6SwIaC95QL8cVHKyUzvQIMy1DzrX6EV4E1JuYWJ
xCNDgXUTJ69VlaoBH3cLxcL7EoqAzWfKrGjfPxIi2nsPodxZvRoDGP0YGS/XGDsb
pQNQcIrrDG7eePlh7XyYSt28gF3X3DlgihHnqnmPErGF9ilhqsu1mz9qAoW/ahcS
qkh8TOyw8bsACRrLZASut1V519WqyV4y0SO4fd6MW9I7wJMXyBU0BrAcJCWxskto
kozxVQDddYAkjsCULvW3NsBHp0dhaGCeQEdaJ81zygegejQXI/Wra5Iy5/rnMQLi
OSRLwCpficanqf9EjyMiUCP/0Z4o4drOMc1lECtNO5Wq5yEGRiTLzfkP+8a//Hgf
CFyX1YJsVLXOnj5LZCbQTNZ8+9n8IJB7mXKJrG2BrbJCexQgq8YmH55s6q+FreOa
2FT1JMWLTP3lK+QL2BdV2Y+lGIW19qm5uv5XBbl2CrHmJcU4KslNW+Ijl01vNtEm
O4oqbrNQ8Ndlwsq7q/XTWjrMX7/jjf4+fOTI3mnBdCgwkB+76FG2SABVWq7fDNPG
UgGKzpA4+saFLdiNr5t/U+91bqK9Wx+Z4yEO978gkXqLtDghEsKwotncmYA69XSr
upBuUp5FhXor6lgaM8lAzEu9zYPYLcuY4JValmiuzYYoQ/HYfkqpIPSxlhrDVNkZ
15v0u0tVqig/d8M+2255cpmo1pYGhU49uRihkDUK6xXJFLukm8RVb2k0mJqbZ/cx
yXzoJgaHowq2LFt74JJ5B2G6CTj7C9j46uxEXB37kDFKa3LD5iRqvaNMDENB81F3
ewoEXjl+re8RAfI8iID+ETUhF9AVFScvc/QHb1QYLtFLBm5Vs3hztECPJ2S3bhFT
AnLd/eKHxrL7WpVPBJ9f9rjI6Y3DdsyiEwHCpw1qWjXCUtkH1T0nfOH90Fy8u2QG
ljfvCQ5BI9aRtn/EH0zXFZNB8GC1oq134yAMHMyY7UkQtswJ/XczcobGMWmy1wUo
+93hdaNEeTkuo21VzMamH+Gi7GQGHu2cyARr1QxT7r6nnnCKgVh5qY2Tw+iXg+nS
KQYgFN4oTtEZFGvvOrAZ7qbzsL53WbjYhwSbVaJaC8ZyI1L0O43cYAREOwzhgRpt
2w5zl02q1sfE9IyZe60HSpsUuYf87AoyfxhezcQRiKZh3jGSuRiXvEBPVZySTjyV
SAsOCet98EIRoWISweRgvWLkipSIePDmVHSMSndM5ZZk3fxzIjKxhHaRS5pFWjl6
m1oCkKJlqVaN8odp49ySh/PF1LQOBzl0Cc+4s6FTjN6HYSRU5YQQU+9RuI97O6bu
EuE8GO6pivEa8gD2aN84BoEqKA9i2IPxjQerAdqzwJ5cPYLqeeH2F5lnlLGdY30+
x0pUhFcEM8dPtkjlmdldc7u99E7SgIcbojEjam5TYgRiXIZEz0D0KJcWzLqu/fZx
+YQBqVZbwVdqvT4MxSjHSb37oZbv6HenKqK9NKzVj82pzaNDq+6GJWbHEtzjlDOr
9MjPfwB/pLK5deo+hpxs5PWwt51eAk8ytX7yLgjf9xlIqW90zyLeIbfglKeeQhH1
sWrl8VgUNKvAR9cRu/WDM49wLIRHqZumaL4Erd05YQmpNt7tAiEuM84SV0lEz6Zx
qlA8DlJAf19skCFvH0MIaziP04ZBIGIIzfCm+4oH070Nn7QPfbfxN9yQ4tCDOjCm
R7hQONPa2bxONJ2BZBYS1CfwGU1E2Q3Sfh8yGYbM+KBaZGZONtw/VugqQdUyg5oa
ujYLgNBK6Njufuon4wABEu4zV8na3oPQ5LkSTwsZhDhWRhHtnfH2N8QEnHZJFd6T
uI3qcV0nSxy28xpAgw6zg4D/yriB6zINOsdWHZavxXZ2s7BCq2G8eshgE44XG/Iv
EgWcvD7vHAbT7NfkLAVLr6uf9X8981LXROSWePC80CirJcm+SeL4NiR9taEmROfS
hu71NBcIuFrLsRLwFGPQ/1UshB+CfgST2eftC0xLS7fejaQAeDS9EKsA7cDJVVNl
NtvvxkX8e9wetE4t+HO1iBiC4fvclHUQNddyNR0rqsdVXqtqTbUXMdSR4JKWnCG6
Z60OZ/5IB2xUEokbsWYakvCuk7ZV/uNmRGiOivtUNKd9/07Xp95kKk1tRpVEBTiW
vBcDv2pWeTNLKsjKrkgQeteKOPWxKwd5xOPyHBwaMiUBxOQtsyq63xDnmEtAt5Zp
cEHbYi5RCH4djR68RzMDiJMC1azFgwK2Od9dcQUPwI7qFAaGuYZ7LJ9R0BX1S9Xw
8VwLH0Dh6qqUjVVvdTOB4stNPHUkr4kQ5WHyS68+gN0TDZBupvJQ0yrn/5KmyBoN
qXBeb48uUBlgcIF4MSU731IHFvB84N6/gNPDuCAcAp1H/A8xjM0Grn9xfBXJr0hn
MWw7c/NDOpy8iKm3PqlltWlZpPyxBUGjlRT25VOp5/Ncbor0+eiL3a4ptoLXQ881
EzHzqdkzt4zD7fVIlcKLIqnc7idAPrnIT2dJ3hLcefdlXrGX3aTwQ3ozpwI3fWy+
kSV+YUTDlu64fH12mMVKiDU7ssLcI8DLrmCmpXxRfOmiKN94V56BKSJ/4IlD8Mhf
nKy5pa14d5xXLzTg+k2pzVL7tO1iN86NycL95/HRM3832i7xakd8VWT8sG5h7h/z
PMnYK5h5EYTfkDpGt514J4jBeXLPG1M7dEzVxedp6uRv5y08x+0onennXkQJ9u+N
1/R9Q8nQiX5ZN64sre2C30BYyXT9UQr4SJbz8tBXRMQc9ZufpdBhS9LXYSTkP9cd
zMk88g+3t6Irx1fSebE3G/jKms/oNaYESk6aj1oO27abC2KqKX7gAyyfHnWxmdVS
FKD3CgMevK/4W1wzWLTyvb39Y342GlX90AgMX+cN2Gz4/iTIdD4MIN+hVNRHjOH+
G25KbuVuP7S12mdHQNdCB4jyX0MrUI8qcPWTCUsqXW7Z8T/YoVIRS2nGm86bgUaf
xYCnZ9X6Diw55MTNd9yk2SVNbvKQ5jZqEQSPmqtJRxazCJDfgMWpryxpiCgsp/B1
mBb11NHBUoL4JsYlBdsuYucLKfK873xqmIQM90SCzGJaXiK+9e70l/fjZDnBsFwE
CqXxZOPCh9+ULT7k2MudXbWPzk0WA/VsADMqArXR3aBBIF+UL47UYsN9puBC4xlT
2IzHCB+8t9IVkxIadmGz++TAQvJm0RSPe40aRulnQIizkzCL3KI1qalL8rbaWYiH
6wqkcKXk9qrwTzOFIHdUgC03aLjNEy9QRIS40aDmnOtkrn007hn0Jb796sr0Rl6r
QilzpaVyP1QMbDGjvGrk0c+gWYWthqp9LYFAkg2lJ3xWpCWk2x5drV0TXomHP2GN
zLI6G0VLWtllAvXpn0iN5dYq4v9VUNoBHQzvviNEPmLOQ0act75GllDta04T0ty+
aqrX9Oxv9sIAO3AR8yop9I52buvgzwf5oHyHDk7mLTPnQZknh/LNllnUee9dI+P1
UkOURm/Ldo8I0jmCcnSCRjMoUsjcNO8Z6QMUIvzQy6XZ9FAh/yqkdwdS09N64uO7
NfNZnHwWhPBNNvfGlM/cM0EuvHa99WoYD8uOdFX3We8H825whMuFxH3RCauucNRK
einpL6v2pEeV29tXo9xsovEPY1vUoir6J3vN8cDSUlKaPjfmBK+w2tMH0IDsUbyB
zhOgKss/jBtW1dyS4CKfZZsCkAG2NXJdX8Il3F4d8URsV80Eq+h4OQcFK8jsain8
5qgLmxF4m1lad6LrEXf4F1K0Dqy6U3zGGfj75Vw80DMWHWg4RRLhhIkuvPJ4yAId
fBUz5Ac/rkZzzUJBcjw2HVrQMfivcPUUJ2DWI/jTxE3WPUCx6fKr8wDDNhpobcmN
jG9LJdwC+lKtFK5loLeE2Lq6/sMgY6C63qTZYMbwEAXjTassXLK0E2F5f2AIwEWn
j8ZGsRQAdx8uw5+/x+ikP5Oa2LTQABwZNwStVs6Uf7ji2jX/LSYP+G6CINuIKo6a
CJlLs2Ths9zINOrIY56D3qVQ0yqSSGQEq1+mwlv9o2phYA7/ml7jCltLgbuMd5FD
qAjkQ6KyACaHSyG02HOcqTS+bVKc+ToFI1hgncR9Aq4kLp+jKVcEsBauGxu+NJFt
ip3Y+0CLq/XnDNAGpYaK/8ikjNKAe2zQZCHu82Csy8jvgPdkZtFnYQJr1VIz2/Sp
MpeFkcs/5mVNgBfipPSfymDHWwNBaUuyWAdoEUIyuJOTyOkJI930I2qg69akORJf
cX9uBkWNtsWMTExrPFohWF4e1VVLtBXh2mowuVpFT91sojQlcNEWEMnwsXW24LNC
ZfOJKzjcHjGHO03kFNndaqOBCJfsOILs0hhnbR3aDWnMd2dKLSzmaSoNMY/AfnEc
14lFB8b4sRjfUoL+xHGMGGasd1/S/O2Kv4fCacpbL2Kmgkvy4yxIOdrm85gPc3se
VeLRxhq6a9g8RyVmageBdYiXUYJkGnn22Ppiq7D3pFnbvvh0o0+nxGCsvv5hakHJ
3/pxozvsQrH5+pE9smBXPHZW/H4K7DdhvpcOOo/vXZfXqQIKefM0QTgld4GUmWGU
IZfBYXxrZh7hfDdfVJ8VyMHytLXGGAnxnCr0l8HlACD12z3VW3ROqCkVXvKRU5cr
b/Rg6owWkANw9UpctMf0KkDOYrY+G/pM+gPJv0E5pBYRZEE5tLdhy7R3mVk4BIMA
R/wDex/Tn2i4oRmRF1LMkIa+uShkAynh0eQQhO1MsJCKOlkZoCrO3QHbfjSYeg81
rg40lee3w12U07GXFALF5mGaXN930G5ikHogppEFRdP1hp9hWorvCb+7xb81FROR
mEof1v+KYkykNijGQIM6xN/7+y2CeXmTF+t92MchAwM2TZQAvjDmga7jyuG0CSmG
GFTz/DM3iU7Lk5wfFGz5aFx3miX//eq4Qt/tLJugBErIY5PwyjOKD4mq8fIMZ0tM
WfDIbSw+1YnllMYD00OxthTcgIoc9dM8wcre2pwhl3WFsytbQosk3AgXbH/PfQbF
xrnEB+mawNV1UExR4cCYlFf/MOgFOjNIiKgZNx9J/vxPgcEHMO+iGfV3jAXxXkJ/
dSCb+gLo5fG/6kb3Dy64df89fFEACft8i4DDPt6MIcUlwLIfzXdG47OKCQexCHry
zve6uXnF7klAx64oHSigP+Na2xXkGo/rUpk+sAq5s0B84CiBPIom4PJvLwlSp3Mi
K4uJRmZA1fgkfucVjtDQIVnNxO3UA637mn+Ys0ib4YdoVrf7wrnts7PIMGmdbFPi
2NnGfom1CvaM66rgmVNqcXFVaZiyT44mQEaMTZAUiFBrCpm9I0QrRBLuOvGPQRSM
E0YiD5JHX0xKmg8n5HBkn5j+SXNymsT1N3aUEDxdPT2WjWfsJVlZUJj9LGtr7m6K
k+osuP48q9uPjHVa59CpmObN9tVKXYkketF2SjxgphtnXOeInjznbvJCUDiaJIq8
TzqrJ/L+jq+oFmpOwmRiJPrGRa78Kfc92NURsB06T/bN/M1zjlKT3YRKTDyYvNpp
bv3/l3rMLFXSMtboDVLm8nwxR2tQtuWFnsYxi2lPX06a35hL1Dvkgl7FospWTa8+
zb4+AdR3tzO7m1w4iuYqaKk/IYNxsY+OjFEORvnx/ARRnbLnHtOkWd8EGECaRKam
gc2eBLD6xncUDrR4iNx8gNigAxd8Lr8q6CknF/HBsaUakjLxBI2ngPRrxbr/HVAP
njuINsb+KwKchTHw7CNWe/1UTc3cYCDbkETaH7yfFcuqJ6RccIf6UNR3OoX9kk6C
WWQeG5qodznT39U75z/pXUCKEmkThWQG/Mv2FDWcSeN82YknjxgqzqxFNqWxKthH
GQU6+btpk3YlW5pZmyvBVwzQtRnUNyNRnr1ugOh1BYtVGXtJd6mlQXdJHhpunbxw
/jr93gmpCwmHnZ/yh7Y1RU5dPoo7ZkSdfShJQzrfFVOos/iLDv56203Ni+T+JRpl
LQ+BfBRRYbBJoObJzV3/Q2N0mGt78Rlf0dDg5XAVPoc1TbpmDc5j3hhho3OszJbO
HjOkYelcEWQsidlPpdGrTHbw59hhjjO9Khe0cAEdnNNE/Yu2+2ifPrE/6Zk/NfF0
a7iNv84zHfUOKud/59XVwycYfWDKD8pEVwznE2ee6rTx0stw1SeCIFNj2gbJ/kQj
mf2XfWv2PjREfwQIzhBU+LJzmbrCnr6owToOvN1BiwJjZ4dzwyDxrmJhrXr/9y+n
CwshglOnCOg1RfYtPpZZobqmOvlc/Lj6BAGVa96hacxiI9TFndZOrGiHLvDAMYiE
JnwjSwhGEx9niqhlc5HrTtIh3aa1Ll/bfsmlJCk9GArd70TfTlvjFFP0DufoeVDw
TfLnRfVvPQLKtqIApfx8lUTdY7MB5/OSho3bfW3oTDsEMNzyUE3d0wbRKNRErsE0
euqg+9CTNJWR9NJEcAWFBAHIqaZ9j+jvXKNVINUqJ4zxJHqmpPIHYdYxY1rnIhg+
xOYOuC5vTxRTOQ39/BmJ0o2ztCgYTwejFrEHFyx7Wi0xd91VRBiE5RGgB/tp9N8n
A4ePi8aV3wdSOiUjJOXNnGNY+/glcaPrMNn07HsH0QaavwwEuYnC1WESoEYOu4qi
tiGCPNXHl3DdnIHhbzIv/j3Ld5t9R1meQIUX4gS17GfOTqiiLInBIJMpuGq4HwGr
dMMdAVb0A088iwaX4AcyQiYg5wey0gy7SB0BESkn4cyfuftETkybU6Zr94KRzkve
4xfy4C3oIsVwCuL26zaE6XGLUZAslFdYL9NVCCRx4vAxFOpuwbp3U6tmNq5JhfCd
z6EAPgx7ISsCCDE0dqfPHB1MlRfdkeXqmPgqKrPHiJNTsG+42vxuhceY3+FzeiWE
PqVueql1ue0DZE/H823Ui/PbmKo1irMLo81gXkTMMXaJfXxmaa8g9yvMuIb1Hdw5
vekdNCDITmetE2zmaoiYOUIx8p+WRh3Ymxgzt4O+6KQXOR+9iEsszxndV8yr7nJu
3NYrmzJKwm7XjcEISyLGJEzD4EW3VJz18wCJ8yONxd+VUvVhx4T7swrRpciHWPu5
1AUMisFmjGUdeLksUPR/Ys93QAkEA21LAMOiTpE9SyxAVtfbQcyNkQngunYi8x+u
8OFAg1CXLJgWqUxZ16RODplI83LepJV5n/TwWrT1X/KLAb26AK4BcD1reYpj+qlu
DdmTfKIiYMGc+C31aebPIauGDsjIR7mC1S6SsHS06Ss7LFcl0i7XIZ/obJpq/rTp
5WuLogf5lM1Tf9yA6UT6hM+9UnD9LSbWLPnwhG2uHuPw1xM3+i2b20F/zTovYpkZ
iQY9s3139fv24o38NjVGjGYJZi+XiQ3VKKiVeMTtxPwEWoxyBu4y5wbh4njIVCaV
3TGi+KJanSUzisLSCAo4aGZxKAPbone4JL23ouoOoocWyoNeGfcbLdCxcZtOAoaQ
pymlhSJwGLZSIBWt0h//qGPXO5AtAdxx2WQY23O0t+s87wH1MhBLTgy2C6q5rMgo
cULp9Y0nHGuCT/8439+ueaND8JROpewLere2kjVkT7QehqzVQO29X2BjkyhI14Fe
lTIUyTbpVWuivNpI4W2FgHQHXdA1y9Ylbda6RMGJArLOvfjcKvFeW4qYstzgaFLQ
cfWoP95+ohRnmep7KvqJpoSUuiHdd3eAXTxV3qhpwTHHicrbLM9UUwYWsFJJOqYn
H2zngzGcRF/ye1+rQFrn7hoSTYIlhPNUW0Qe0Kg0mKzFVkllTamvjMGFrXQJ/sIQ
Faxxwe4Ez4uvdN3Nj8lUndUtBnESXjUWJLJCjeYUROg/Cgx0PRHmccmzFsIGVmBB
Y3mND2BsvhTtAtKj6csyN+n8S8mjf6XiVTfOXkwPKEh0sPws+yMWgCwRWydQPBVR
H++0erwwEGniGekO51Yzarc/8bAKsVeb00H6TtRKmm+L0uy95x0aCET9ACuHHSB3
PDAyLx6UeVDsOmn9GJSGwa6skfAasnogyP6CzphaJeQ7MPyLCPYnVWdqSnIcCEBT
cY+VozArV02Lpgx8vSzibZu+4TlT4syFP084FStZMeAu+RfKq2yx+QJr2I8rTXSR
rb7Pury14JM77uUPy7opHtNdxHFZRttCR7jeSveIxiq3mgfvUB9efhlEBHLLnxD7
3k+kTGSTL/SH/ws2sLDniEHcnhrTLqt2oOu9m6zmbSKqFujLO8AvLlEKk4NjVlv1
+hLxyl4A2mYCuCcWHBaiXlg8tHYCiky2MgWfWuEUCkZ3iuAs9M0ZBamaZglsVv8y
v2Z4rJiP/CFySQodRGUdbA9fxAwzrwKPB2SKvhQBW0GYDeE6zQ+MiBTobpcRbfqB
W+QQFQLrUHkMdyxdB4hpuccIeNb49lSpAhfcj3VpaOs7fUbR2fd43iV9hsTbC7U6
oZZ5vpRRxugAu86Zh+fB56INEWiQQpYw0+LV3Py2sM0i0XxqAn8utaIrfGu+pQNl
2PQaPQOwzCUp273uB6FrL1NV7YuXjjOfsFjy8yw8Q+ZIV+h9VQu4OP2cbCYxAUk1
MaHmUsJMlK/IiU5wr9ooQcjXHwKVu74myU+pqsY6fDkqOiWZrU1xzHreUCqDycvk
PhBTUTyH1dlvZMUX/Sa1brsH3y2XKPxhhsA4o99AlWV3ERLRlyftLM9kgMVQaeh+
s7gzyrPtWDbluiOVE5PMudtdFsiaEiLVrywpZK4Smx06dhfpbkeh+NPbS/lOsfNA
+Z7uQXfpA1O5zfSetMg5m2Pdk59oRTLvFoSNtCJp/0zDMo0VNdYH4MjVcHLb+yA9
WuzMYpJ9wAXpKtmbUnGzPfv/mP9KylVS8xCgs3UeahChyeRzZarj8ihgCXqAH49r
SQvKtNyy7MmLgm1cHv9w4uD12gxCUvLroQepvDqct6Q2g6aLduO5z4DGUUmPyMgs
rgWKWqJb1hEDKSeLqjZ6UxAvG7zHGn5A8yC6IBer/vhOvhQGEO54/rPyzPEP5UuP
6kTb+hNq/NutoAnOWA/ZG+WqcAFOalw03uzEbtuoCXrAgcv6xF3DigVsXYEkWi8O
/H5r7HRY1kwqRPMF+zsaDJgYFQYpXTUHYPld6uTWHCE7OhkoXM3MWuKEvlHHtPbE
CZn5+o7Vvo9jFLfO/LMOeOOnbpQe0GRoaazai1JmPiUZRFOFxDE8kced2BkOptgt
Djyd8qORaPCvi9IAy8+Yu7HVy9b/X0aCLXtdXT2bUxEdFC1C1aTYjQsgpNTCYF9C
Ov/YoYNlfhn95x9dLn0uVVT35T3B1BylKttioD2CxZk9E2scEqeBst0pTifcbvUl
iuugDHfcEC6JsGDPsew77X57N1gJfUFtYxsKRZYUwZPRwF9Icpy1kjQ5PC3Sxauw
2V1tJW4AB5NF/W5A6UHm4LbVcO1RA9kqXXa4Q1ilnhXeTi+HH08gwePN8dtPA0fb
9E1aWNCTN2Y8U87TrpHbaazHy8bZehf5b8DT+3chNZ6g1cEpkWbumZx7OvA+06K3
ftCdfLM0F56U2ibZOj3Zew7YQb+/044NNrlC23ep8dONgIMC+YP2hj/ZH4p+mMoA
2dNtgYWEE5zaB/4qFq27GaUF80jWzFnofYy76Jlb68iOjIpDoXlYMWF57Npis4Tz
KlFCkFAsjwDJQ1pbWBXx0eckou7+MlPre9zk1KFLYQdoCM10x81jTyJ2k+jHYFuc
Xe4eJlgKnvzx9l9mBl8zNmEPDzqRcnHKGsUrqhWosdu9aOQlswVD/BOwKo1I5xWs
kQ3KN7PThZ88NpqAwDhpRmqMialnVahowcBothb438a7B2/v/+hGCC5aI36D/RdQ
0sqdHarfIdnwzqYgzxBsTHyHB2wuY5VgjfLaGwG3/aOUO5RaHERLTbH934WW27Xh
wg+/4fB9gM2F9Qmt77RZk1h916bescWq8vZHRNy5CSUvvz3pBW1QEES7gLp8n2qG
FKGvhK/44wg3Zov6BlLK6un9ayHfk0WLN1W0Q5PRPFA+KS6Mqbdg1Nvpr0L91wHs
eoAGfzftQ0DgiixFdqU9qPguOtVeu3mOsBy+z/h4aRpyxZNg9LUp3jqq8yq66CKe
3Rk8pEdGFRK+/YWd5aIcbiIVv/Qn5dqxpUK5EHi3+/1vpUlfamD7iqXBw+YKz1Ao
WcpKtli/xTSeA0A3aXhjqYB+w1Xiee2rCaFHcIGxFWDQppuy3lyJe7wuXhPkG/d/
rUhUvs3P2jGD0BdxAjAaPA+EjiUTJmSd32ID6PqRmJroet9Tdvgl7Vu8SLaUmU/1
vK6cK3dZrkzJrXh9v8sBeoex+LnMZEIqa6rXz7VGapJTxfB9BX4kE+luMm/im4JR
5PCPHDOJ4em8tsTX5C4/gnHPLRruAz2REc4FJD7bDGyVBGgjDRAJ0ipT9X6gPIwS
TF6axoS0RdRoNH9nwrUvrABIAo0op5418ENih7nxlMEv4LqewXKCJfR/XEoKA7B5
Vm0GAwRVwPalKDAfdtOFrD2zYu0Zi+wUKP0WTUh4/S5i0YG+r5QzHndcFV3Mf9ll
LmS3tA9kTFA2eCebMAstybK9VRN+T3VCJfa/H7uktWbySX2ZtSiPRSYFM0BADYBA
nr7AuAgtrcXUFwMEI86tAU+hz3nw4+MC8C749RBS7ZqBhYPRWkWXZbSSzw3NOwAj
EPQN4m5hpMUELBqExA6IS4i2ylqyu/0YKpGAqjrRxCZxy7KB9BidSQM7uMVIO7gc
/cwD6fZqyoWwjF1HJlhjehtahIBraVj4HG3tRHdo0QlOIp9bvMZvPpV2AlAQbGhY
fETEA8t41YpGV0j40izwiqt7O4BGB538PNJO2H5ZA9ofMgzbqlx4MxBwEg0qW5uf
xhZlDUSJe+UR5NliduDzM9SBoHRloTcmswAJvI5cC6/WlCb8thV4wLCeKDQs8DYh
ZASl0XvUjfoRCdowkrqM9RDqoutfgMPOHaUqbKVP/4QiI8pzb1mSsiJqdCikNFDq
m4B0Cpnak1PZPffcj8Q9TfuAjGZzL41etJ4sI4j4LPC4rFpsx25dofrbSkKmS43D
0zByqgonlprUt+sUQjb2X3YRT+MpjeZ79MZe+hKGLXevKdwax/TQtXYZtDSNGaWS
tMOe+qxcqJ/BAAwEkCNY/lqI5j0iFNYVF30D5CbVljPqL3XowxUDsYghpRW3op/E
FGL/vZXcn9Vo8J2iCHZjLs+wrpGRsNJjJ+SBdCP/ShCQ6uaI7JSAIQ8ysbcX+nBr
yjp1MN6szzCFh1ZnXWPd3Gxm/Vck0D2DgcAo57K4vXE5rZhOjnrKun4bNeZFnRk/
w6sWh5w2lxQs1Bp8wcobjkoZw6sYQR99nmbtnSlyA1i+2zCfytlccw3lW50l4WEy
w2BPjVCj9ajy2EThhTqXYGlOMeK8ACMns6CMGWA+GjaAFVSEANN1+qP0eDklXzNq
Dz+ZszmJREgDM+YhfYRI+mkrxxhkYz4xuJHIKWnTEKkVlXU4uMF6u/tI5m3cyomI
IMvPhUWHknfmbl1K0ucYczqIm0nTKMhEAGJ/ag5ZBG4cl6K0PqfSNvb/fSfyqr8e
Dm+4W8+AYa5RjdgxDxv+Xf6GYf/eSjv8CXxTL9V2LFgVaYUesx9tuxYfPeLo2ryx
N7kEziFJqwLMSUkL/GCdlZbem6OSkW/V/4GX1biNVt1+7USbjEliLwvSZ6H+9qJC
D0E4FU2XcVc9zb/f6CjMLpXatz1ECf4in8wxxB5YB8MNJ/c/dORL4a7aqH4is3ew
XteUZJUQIvOORbU9vu9uDSpmabbQr1lHB8y65eeipJoUQ0Od8ITGRTpVFWQ8WcT9
7IM7F3bwPxCIMOSTv8W1dtD8DJ0XnODXDHIu+qOz9Rcl2lBrZ5efZGD1O4ZSTu7t
gCsd/X+nrE/x3myCsQc9KvCyJDFjM3EOFRcXDVEy86VMn95bRemBi44PeL5bLSV9
5Y/rak5ogj63QlLWcNt1nmh3QbhxqlobFdfrQs4WBz20CXuIpI0+ldg2ko4X5wdJ
ljsd6Yruwp/Tq+tyGRhZeiih9QZ9Cs3ccczMrF3ctl0TEFUWMBpeTaO/Jq7ML7Y5
taKCXHHOZXulcYCnqdgqDgL5WtAcfdzuB0RoqjWOZJrhXWzfov5E9HcIxKqHHUzs
H2pXo5hGDbJBbSMuxgIa+2my/IGBTZay1z+jY5ug7wkUKJmegl8qXIm/sHUNsbBi
KahUfIsvslyuezpLh88N62BVbV8s5u4apQpgIkl0ZH4wvUUinkjpnR0/FfAy/2Sh
fe+i8xXeyXPmn1wyjYUAtX966oMaTLeN1s9QIIkbjRksxw72RiXfrApweaX3TpBZ
VsLW+cpStO8oCVvNDnGGt5pvEFpxuPi+VLOa8R7ZYFqW9NhGHVl5gK1Q02m9j3hu
rNQfFOHTR2df3dkYFw4IuzRzHpOkWJicBs2l63bnoaS6ZJpaI3Ac2gz5rlDk+JEc
CLqXbZukPik+hdf5Owb2q9WEXOa2284QTBu5Rwp9XuPhSSAyciAadH2keBVL89cq
r+8Cwxw15IgJjCAYy8HsMzmJFrotOUxkuczw8K3/Lc7aOpbi9EKlKOoR1yIE0gG6
hAO3CSFMcyQR7L3P8nYjbDJ5YVhrOUGkrr/5tavz+9sBdinlNGveywPerlOfinun
GLIfZbg3yWNhjueTPkB0Q+8+92mZ5lKK2v3hYj8d0tXeEGSepO1vmSx67/tNQmzx
gFMmp6xV3eBnXjl9icz7scLj2Xm5J5qXrc7pSEYqBMNnhTJwMatOzx4vLpQlcgRR
NEaM1p58sjSYIo35wWyhjW90wS7A5vWL5Hlge2fakJwYhCW/dZcYZgqUvo1Vj6Mc
ME2LX370G57xXD6voXv3T/xBb4eK/jZPVLTTddISaObpg9J/7j+LakzaGkG5eVIS
9OX/rKpIMyqfleE7qA4mRvp0UCiLWiUUyz6HDblofi6BzeRrgLpH2rzMJlnyRaJF
RkzDs0TuRHDeMGZhSEO99kw3mdq4UmxBbXwkL0Rof+sTbaXthFxFWQ3JT2jQg/Te
RgWHiq/Z8ZoeFI7Uf0zW3zKDAMJlNy8aSDjo4YJQSo3r0vb96sEA3tostisEByuR
DRh3sBIwUnUWZOn1H8KOcCqB9LSfpXK+Nck1/geISsQ/kyh8Zm1KG/hEulqOMYcm
JtnjM7f/qXB2VNNFPmFBug7hC79QJXTk3hQtyMf+2h8tB/l+AMKi/yDYwCWbsCFa
kGj2Q2uUCcO8bTD/LEDtozy8EdaLzj//Dtwpy8hk32ey3n4LYz5G7VxzuL4g/8xr
AozzKykaygNpZpWufbPtikN0B1lDODcew2sc1ovozPkKRvItXjvX/tGoJW/cO6PC
IzyINrXP6BpERV/40Ce+w7RJVn8RlsIHM/P63BhC/s2t1hkFv7rk2SoF4wHrds22
1bFhmQfAvRBp/llw7WS5d5KH/g3RT0HsxYgtVrvXzdjvo1MLncoxMMMyEvZuzAvt
QrVa6Qmn3FxzA4205dJrP7s7UmVsL3qF3HwRzYUwgqQHZTEnSRY2X1B7JhqWCJau
7DWuTFwKa5VFn5CMCCydHHE5k731hxQiRklWZn1/rF96delbREPK0N8EdpJk44ph
FdqyWvwVhDXdabGgwMlGUdiS/M8bt8gaI/vw8nwelwwOTMmMx94GVq/y3BqouwDP
yZJB76YeZnkWNUbqIj9ZWNSgBqh+xXtcB4lBgMP8qz8HtjBj+VXbQKgY/L52RHwX
mJmGHYRJi1VAYJ3sN/+D7f2OuKSi2pa16jKRIuirtaEtweAeVhu05bj0oSyGvIYI
qcMtq3aDW2K90rDP7pSTSTL4VR9c3iCfbagZawoLyO2iyH97srOtg3PwOV0UruPL
D89yylXBeQ9rY4XNoSRpL4bENdEsPYllybsft67j02Oy29kGE25t/sO99IO6Ui41
PTk41OmVIxD5auzMYSWYeKAfHNbaOiNhQDZ+aNfexzcDPI/aWHtWqrBHduYs5QJN
QgW5ZwxHv/Y4H2ttfhdBJZWQ0hUW1WkVGuVHWdtn0Un+6xJsN+vks1iD/Hq04OlG
WlaBKjNMbBU/1EBEEMQQTOeiWxrshzjgwFoIopQIGfj1C5771ahKZdOYlaXnVP6D
jkIe/Qb6rgDj4Cx0KKDFiQPFD4NY5TFZLuFTG/pel3IsL/QtvWHxFK4tMTH3eiqV
eZH1pxUOEpK7Tgp+spGS/kR2IsOC7eP5x2ZiSLEBB0tCZ4+HpC/zwR9asraQ4Vsf
SWxSgW8EqCyeiYzfpQzK35MnFpAuicDRIs/KbpY1vDzvH/Rsow8i+oYhktEcLa8f
gLUIhkFBpkXeuwUkWvKoGQ9Hrmn9epYfBDCliUqrA7xl+p07VOT6ECUMcq4x8zuB
YnHlw3AqELfxnbbohJTOFVqZH0Rbgv88O/3QHOhuQF7YQhRxQIstUCDbbfkGoLDi
ticQS2UDyKJJ6ZRkIJ8dYXNm2L8gXUDGJ3ceo1jgIhL8DipYepNggsLDoi4CizjH
uS/5p/FjR3LXukRg8pS9WZ2XgdeHRdxbvjT4/z1u+3/FyA7AZZhuBapZffJ3GGB2
fBHlmgb9usOnVVgCT/W88zpQ5vPBEq/+wYAngw++Jz6nl0ZV+rePZlTtr/gi/SJJ
TGur5121sCpgy1a7OIbpcE9v70rXVmVjZHoUR5yd5ZhqLzSuM/CIRwLVBmqlqPXw
wKGCd7xLjoA0VWxdbdQEhujCOXB596Xw1RTcq2rR7je5AGskQXa1+8gOheBG6j5o
A1HMynt+6nT3uaxeBVlTEqnQvTJM8Xd1iqcuxFP65NIf0RScZfUKHgiwOrl0JD+s
BtNC9ZwqcweTArob+gHP3weNvi0p4xiDpRs4nI9r1PuTiIhlF0ysu6GxZ5YrHY9o
sC3deKuKOFSxxKY0ftO/j9xsdWBg0RnoB8aETbzmOdRGVo2L3tdvKnvQFEVhfM30
NDv8qwcu+jF5XskoqBNB5KKphhpxk2jFN6f7+/INpR9bCVR3NxNYxHkklO1D3/dN
FG3yswmRSz6VMg3P2++lvVq2+2Wr0Ng6a+hKBFpemzsNJSZfyjqZ0e5lmCKo4nD/
Fmnuup85O3o6Vz1wpx5jX2qNyXG9Omrey9065viB+x+H5ITK5mmiLqzccbytyj2W
cRxgudzzSy6V/U19r1hUkP9GsIMXqP7KExcQSi3+Je+NZqnPmwQ/Oym51J54WwCR
SW9QGVAmgdDwXVf+18Lt4bI8A0cX8ZuWoq6WruQePUk5EUdm9np9gjeNxZDOGK2V
1jdnzfNzA17UlMyePSuBNhGLV7wvLDFZQCwskX3AoSqIVluz8nnFPYvUbjNOxc9f
m9GiF9bLc4hnU80g8f2M+BqYmDjng8AzVRvjSyEhfI25r41QyHTKV6nsZLheuV1S
0ndQ3OJL8ZR5oIXcK0rZa55Tpc+L5hDU+zfKmgifnbNADBAGXpTDHwYmJ5D4S4tJ
ILLi/MLhHfH4OB5lCExZSdAn2RKPYB0fbMWAs17o4wPcNgWs/5tigGY8ya4NIqAE
2bEgM1WUfxCNr4c+P6dnH8gExLTDE9wGO/HnNP8PgxrHWOgg9PLcTGXA+FG81WDY
UszDywSH+WnIY+AUSIv36EtKAadkKOOGtwPKP3bWPB2I1PlbXR/ZFtvK8VAvlCuT
k6cWD5Y53i+BjCs+ozTfC749nJkYM/+TbpyGZhtZOeEci74vr74N/qz2wcOFUrPa
oJ3IdV0s6S0aSKmo6XuYrRvWh2l9yHUtuep/z0dSuX1xUQAV4twQJHbQnsmDAVVW
WKFdrI253Letm1N1/9AIbxPwNXYpE2hA1NVenvMOUU5asDa1JKNlAAbNtN2gDuC2
JChckVlnANzEEFer3CsV5g2eIAA572KdQVl4TPGqZ99KRK9Mj6NdfwFcn/VMkKaj
GqIWnThefK4w7gU4OoDn0qhBFpNXjwYUlnmizEixEmX9Te0nMYGeF/SvcmPWOvNU
tQHWTuij6/Cqh1A15fScxas0vVJGtfq29/FD4V2ME6tdhygRZ09fOct5DWm2ZTRY
fOTzhIUOkMISollLOgHQkmZBYHFGT7XFY3upAWUqoozLuew1uZxbN+qM8fI/ULfH
jNvU2e1yizVI4vWwTKsVwO4M/8cYDUq3fCQezPn84wF+PO4kJZcYkgCef/YAPaRh
iZyaJfb1rJ5mmWKbgm+KYUGQ+l/xo3UkPox6gvcgsBdnrRS0hggURXv/Kxbov3vh
hxwS/xTOapVKTg831ZpHItGqTCcrIiXKN91PoPfGLubyX0xyM0KEzsk7Y5cGc+TP
1ShgNe/zhAj5swz/ExZA7e0OYiDPJ2rpGro1caCxn6b033xWjmIKkxUk1f5OSnSA
WLt3e3f+J0O9Wb4qmTQOBhXfxPiGQrrhErV5nqvCw7HorYEZmHIOM6AODoiCzLGZ
mfmWLbdls4kB+g81CLuZpoY8+86pZIlvtWRccIwpVZmP6Osaq3lICj64X7yopElB
KBxUUEd5c8JZv3biFhzD4s+z3qkxMzT6swQEaklMMh0cohcdcnAwYXV4PFqQnKSV
oM2YBXH4sg2UzIR9WYh3113X3IhxQ0rnEPYuwos7OUfBuLXA2dq9euymHwYN6d6V
D2BFr+ky7YRzijpw08GXg1cAQrUuy9zWpzlc5P+GzTvun2QhatgtYcB3bRqIqIHk
L/TzVBCBa+E2pC63xBOWoiz0StUbDHiNZlnn7TuoEw60mLWtXFVdskY1i1WJqkqs
kB6wFAy1ScZ3IDOE6lMrsncyGnyFxsCkbblkiyBTsS00vnOEw+8OqjNDgtV6rmXn
7htp7UUa+/DKxE1gPcCOcUzLUnCr8aY+oKj73SUWc3yXioE2nXxwEn+SM+kEmo5F
/LAsR4aWWn0rNkZtQGJQzdsT9sBxDUCgnWJOLRjur0TrTRGF8cELORIPZbdXUTPx
0qtSVPxwF8UErmX8xRwgg/rsWd/iX6REKp05or+bvBMrLNui6XSAVYqQ6+qAr2gD
wzxfY1rmaue1iosw1S8VuSUUWrN6dtISR7ixpgYCwRtxKIcCbCjoiWovtHcSjKoL
yRXzxq3pkSzvO+MbjowYhFAs3gNec5kmcEOMxyp7GpsCczw8fa8L6Rdk89DXduu7
eyPQOMesans6A06SJZUTqRtTmPuSM1dHCg1nyr12DvM4h3YpPIe2e2Rqqg6zzSl2
wqEXHg32tqyUCW08b65IIMF7T0tKyOU+/G/HWBIBZUCIE55iK188YX1aHsCAZhyZ
z0XOKsYe4/FTnSU4jM6vD7M04fNT07SFDi+uPPEtKrTB4dJi1UcUn3T/s5OfzXUm
FECV3l+ElEy77zAeuDFppjmPjMSmTsRphxTd5QC0ojAskicPtP2wObnDDRVL/pnA
V3FMZe9VTY+f49bJyfSQUHks+reNhsRx2ORGFt72siK1SowhPf2DeYaUPJVT9ZE3
jNh882TDMHsKPFCAt9IBz0FsMl4s5PgFUiWFFheIg3EGLuhPDJL7RXQApahpNJxX
ECvtKaSLNuHboM84qDhH2Lsj+Fw09C1wDJNIU0qu8+wuHQnhULNGcLj3bjkIpV7d
VhRRWumxap5+ytUICL2TnA9geqn+9MGVhDrvWIZN88NFXbdaQfHD8Pk79BRCdtZH
vS5URpjXWH4atZZA37XNfiQJ0NvAiPYW0cy+/78GEQvrdmJtp/w4OfqVpWMbq+PW
ffjDcFrO+op8qgPgLQs4aGJLEoFbF42C0NivHhZ+9qe9k589lh3cBmHhpI9lI686
XZdjgTEkcSQVnzsdQucv/8lD7ShiBAKOcKf3mEMuHg/nbbkdZi2c+dpWajHyfuMc
l9zOuq+2LNleIRECjh0Tywcol6+eeu/xouhrPtAj67gBBaw2IEMI00zDCc/60tIy
l8XgecEGamSh04zz8EUumgiRGfHccFiqmwUfNdZ24GKhoE+jRvZfqRjs2tuto4zx
l1/yD9YRniThq/7lZUzLFywiiaApBCvMz7m+cjkYQp7o2cUr91ZApgASCkp7KIV1
mNS7cde74HCglwGvB4LnWO0tQiMK2oMpQyhZX6zEDCgEOAqEFtdhYpl6gJl+KAxI
pHflev+V7uFqD+uo0w+BpwEfzH5Om3igE1VxGdJcfMrr+/ZcjoFYyaTgnDi2uEAq
yZiHLZFfD1zwdzioHU6MSsisRUKhQmwI07nTHkqnEj5Rkq5ruitM3opbjIghA8L8
sAy68UUNBFDmPhYa7+k14Lcpf5B+k34zE+O8RFACZelUyS8Fwvug3o0Os28d2d8v
H3vA3XfGIWXMVSxI+olghuTGAeAxhV2hI3ed0/wqBM7kRIbn0BoLFcRYcIot+2Wa
O8e6C+BH2Tx2KqDCHscjPETduf4Cgev2phQqTVDG9p6o2JHhRZAWMhs28+Sl5XSt
rgGDcf6RJNuyP5OC3WNuKyHUeieKyHlGgIusATIwWpq7DibpFm1OKVRiOrJSGy0k
fwUX/MryMR+CnEadwu0KJ0vp8k8pi8zgXSqD3/QIxfmeIUlzc7VEzU9PF+wuGJJ5
EsgGcG4G9ZGAjiuow4tlhZcE5sBZcbVJeyBTkRy/Q3LXCS0f7Y5B87OTPoNHbXE3
vQgADDjf/dTVWm/i6YA2xCgjUvCvc9LSCpHvbJgPea/ykTFJEGcFG8MmKy1Sktf+
5zUrdBHoSrQKLTWkue8YndGF1UBb+3H+pLxM7ugDNAn9kuPj79TMMpvOJdfOe9NK
XJUFSOTHCg+gpg9IoGpCfV/ZJ4HOBAXGjxGhyDo3xw0h0u0eI3bw8ojw8S/royK1
TRYbREExMTFaeBOLWhw9djxfGtf6/jscsX/Bh7yIwXWeaGcfs8s823fiToYc/aFE
vGnzQVTvUnOD+GZG+Jg/4RY2iR8oBVHq29+m/RNp64KXFBnbghGA1JgXC3QQGeJC
8eD14FQnnKK59wTQ2OUi5fLloCE+m+umOF5Os+LdOSMQVjgLoDWcKuFPZ8KtIVUr
iT9F60rPGE2tOE3XkeYs5+F6cQPttNRzf4yDrP/bvzwvjiyPfpejd5pPhAHCXxXR
e0R2mZ9oeDaYzjJYAypyVGnP2fxX1/g35l7//IvHN6osxKJ0zR2muALaH+EK+nPz
m8mJn8IdXTlRTdSoke493vB58UwYbKng7Laz7xBRrrTZ3OuwSUw+dVv1eOjQ7dCs
LCHhCq8SCH2gAUtJ1bJxqQRvE+dSlZ0hPAVshcDH52X3RlQh1G/vkA5BAQOq61ap
EY9Nk/2HCpz6DzqwJal6BkAcPK3mAd8o55KRLpOUPbTHPgQocNi+uD5RILy9GztX
XWt+qgAHgZvQx39sCAcYtwbMmFmgwinYnaSNy3MI+EYV4x2PEKhhuP9T6lr4q5ya
TxVd5jIQ2aBvsyb7nFvyf0/ttyKjmkTrlNH2oE6C8SyrzJb5iGf6Xy0LGNNq/uIX
75YIcPv8rNXQOlcObkLRTGb1SO6bqpnEsZCh7T8lsxZ9x5TSFFy4uoF+vxaYvFDQ
hBHt+bQzBxelcRXsQ79LIFx+yTOGzjRGoLmeM9P4zQEZSY729WCXwbYmKw0TTRvV
u0huR+HnZZxl2JMgYrjVwbJfWYCvGMU1vq+Lm2GXpO4leI0JVJ9W8yhLleJvjSGP
6LaG2D3k0otk2EDyQh4bdG0JZI/UpStbqby7XGe0CZ7P/F4d9LrBBx9yx3crhK4E
zBZFWcoyKdPf7NkZuVH5hxB4Y3VknM35Bfaka/lNLtv59ishNwkFBMsw39mXuD6+
BTvwC0i7gWnGpIEqk4NEEcJK9Q3XM88ny+Ibt48fJTuFvHqzJVk15XwrjN5yJct2
bvcP6+/WWSguzBAsMKUhf/qjqdM6K8cXvyLhpkf0UnUR7KDLVyzvU32fZu1kM3Br
Y08cy8o9uzKSDxzPQRlRNgtSFa0ybyfXF+XSVO0TZpin0F069QyccRtDQ3fG11qS
koNu5qpiATa7CFGobiYpLGR7nXOIc0k89eBKyEkdsX8J+f5tNUpoeEcFTgaQhN4t
HI0I+IHH/a7bdsrVOlNWfKrMiNZUHPRI44ki0dS63Gx9gL5PM4xahFZNMdmTZKOS
aDpSx1baiAgH4fmZrMR+sPNZWL6ZTtP0JCP727rPL7f9rquv70R8x01UVAeaq/tm
fq4ICE9h0Lr9o+F2YHuDQbgEB65BqHBeEQQK/SYQqsRmcQOSyFY8Gey3bWozN+qq
JYPBEE21WGFyF7rt2P6l9NU8+RLwSsMz/5GDXnn5u3Ia+J/0bQTIOhYL8YRpuUc6
4pi7yn4le+IBJpXSRtDoY49wY/4baZ7EZOV/SAswHjji5Lzw8Od6Jhlqng1W3k4o
wyNkCZNWsgBFnr+pqh9jMwhbtMhx5tYDK/H/L1T8/QrFKQKrhINzpYeVKcLWhfFO
8xSVEqyWdBKbrRtYOjnLn7Ppf0vXw9235RjxPLa9IVHozGI1F1FRgKxh15w7Xpzc
qBwxoT+qo/PalyPmzAOgqwZcY/qw8wXTCZgnvxSXfAETD/mWSX0ek76xXspISQL6
vpB9ppapH9i2gXWO9idxYPcRH+26LZHDoWqaEBlHUsU6dh6i9FnpXm29+D1ksEVv
MQ0HhqGdevdiz/DlaCLdYOHlWPu1m6UqfzlJ2k+Rx5GIYDzH5CAFnirxfWf3BWRM
1pmD5WoPC+4Rri3lMCU/rcXUz3x1mcCpyZYX9fK6+57eaZy31FCxoX5UHtLNQUOZ
SY10oXi+qvYYUceQuD4CMIAb/Fr81kWOTgB1EjEp2SwHfBpUPg7iEvFAOgOwBHRh
CMH2nZSnaHfdD+qFd3u5uUNsy+/Y8JBEjs01AwTolv7Fx0JPW+F4QYBJzk2rfxXJ
eqeCIPD9SUUCFlyvUzfGaupHSmFhFyG0R7ROLO11u+o5qRqkhFeo0/x6cYeRUVaA
J0ESDLzo/nzcQnoSHLIxYsYyhRHIWHoCsSe8LkvRLiYYOaJdIpbOjXNWQCwVqWnt
pJinUlG11a1na95TpPGSABIYCwC9pEvd/wxv2AfZjebxC90tHCXW3sqJk/L7xIqe
swmTPO0M9lb+EZQXEi02JzG1ZBk/REDpuDZgx0ZTRjS/zj+xN1P7XxvnkV2qcc3h
B3YuY/aoj1oN6vJu+olgker4c0ll48RvB1an8HM+mqu8M2gihBPqluR2o6ob5dlZ
LDP1SxSj2mKPKxUUAZde140lUaqHJ9Fh4KJ31WksEHZHH6Mx661x/bMwPaBXJkCM
X3gHjMWvtbCM0D4HPsv/J4a0UrZ1kmAOP6pCWzVlfqZPHsM2K36Rre1gUnxZL+Ou
TVIcTujZ62t5PB6m2r+u8DsPIzyBPPMv/JkGTfXQVtzUr5wrtPUziyccvGLo93Na
L0RtRjwkt2Rl7N0+tu4SB83Zo3Tyv/UWcjzOqpQZOTA7edno51u/NSHZjbmT4Mfi
mb8wIr99/rxcGTGuguGT/OXjE00gz7eT6sy2tN8K02s0YfCo2OIzCbb0ifbyQuNX
0AGd6C8J2B211GoWqPKjmqvz8C0+uY5QGRHlo20dh5hKdOTnEEdnRlkcSR4wRjVZ
dAu1GjnwgwSlBR1t68h0B4vwQmKl9x+NDrH9PCOE0zJsnzB0rQEXz0RLbMFHilbS
FVXlqA8lb96+6rFAma2GX2vwuqj0C7bfgeP73tt+uE/jPNodrCMk63WITNDR3UFu
wxqQe8I5JGq1cD5JmBygolN/dV7HDM34UjkRORAE5X78mmfPRpOwB6khJDWRJzAC
PklbG8p1UBF9FgLwNe5RziRdI5co+ciSGGRgm62RO8D4dCg2KJOeBYfYpLdzkUuf
KPM7v2YpOr8ObsnzFX7Rb5b9KI0ryvf4wsfcLXag4DgUJe40cjXwLt5yCPWOD/Dj
6z9nPb6LqRSCF4U8p+eo7jSdg9w2Rvia9peLVX9ArukEkMX9dgUZ7EZnP+JtljC6
XtQme7YU1HMXgcCmohe7zOfUEjAOhKUkZ4dV0EAasMiN2ai000JoV8MYbVCmpTQ2
P65eP6FMO3NRcXaDTtm2H35hcQj5lJVq4HIDL6wFcAeaO9v7AtSBJexVPOifcDEN
iYPeMz1ebYpMqZ0GSLZ9eIHTdR4uy/NfxX7rLyJ+cvO05dXY+SQjQNyD3A3x9fqA
TVQHpIzkbMordrGh0MUUYHyQZ9VLlUYJBLtenOt6inn5OvJ0BUbQNg0rXbzvCI92
n9p/Acni3JcPny88/NNOIPtJRzzOe1KKSvvcGO6FKRPTPGRKqjuY/BnWKul71rO4
PfL2cbYVr4s+eLod9fYDIrK9d7ezY9SdShR0B783KxjVsjqlOh2wsKdwn1Nq9Y/e
FQ5fVCWkes1IClZ2vJhIfNSFTCWXht6QQ7OVLIUo1aDwjTJINMT4zxn1/tJlTT0S
1/NWnlrAUdxTaziwKCF/SKf/LVMAohwmEEVioXuInKUVUsvhrAxgHdAITN56wtY1
Ew3romWdv9D5F0XkSFhYSSpDVu1TOqUcJwWEEZ7iiLVLihKfPEICv27hVooH3Kxp
9COSp0KHRZyHlNuJBHATCkPfLmbw7gZ+1CZM/beHXp2jPmvnVplBtaV72c3v2L3/
whomgG+kUTnH8w9RbU3J5NC43p1bmJ6/6lmCDLORPeViUON7E6Tva/gWd2sIReAG
8QoPf9zrrGOjU14ZUUlkb7pMMW5OIzbUlW6C09hxOhE5c/kVQCRoOEXPLEZ0BKbx
IMIydzYAEObuhfNZlcx3b47GwKsA7pQSakyrdIq5gbJeUrRBYjobgwVIdwZqroEO
UerWkURsv2LitOop2VDiJadCkedPzuBbwH0ikvFtrolyNw2TZOJsHFjOVGRefGtt
vLLrrkkyOGtUzh/3cuYIQ4T/zLjJ07wM3vcu5GRJVT5HSU/Owynsga4fRqVwHpYW
P1JBSrJcW72Qh5TER5qGeOp9AfEbAy8L0yBVHq0hWa5NVTR/np+8UOAl77NYbUNq
1LfOSQCOYtXgreh9Y7bjAHDXlb6cX+rMDM6eYsl0OfZA+jw7YVDDl1hESdKu75/J
cuzwCUdC5nPAiA/Uunvf+q/c2EgysaDbwjba6sHvTrky9oiWyWqkdmSUMmaszgfb
PoPtFh9dFe/SoOgkGOCjYYDxWOVJm8h/vcaGT/VEwjIHpuVnz2Y6nN2OkgnzOBrN
vQzQYQj+EjbhL3a0bCueyelzghlX1vNoHDdyZgDF3sGd5L63leS9AiHkmFpaNs29
jwPEoK/X48hz1aSU+6jcOIsx9QnLKfegYjNLT+w4AjId74/UEoxWHpmaPWvhqGB6
tUSqlx+D6jTe42CQeMnRU7Z0XorTAfu5fyMtmRTjVjwowV0OH9eESDJ7pGbAqxHT
Z7b8P0IP94naAAhfSnIFWAHAwJvRXaALg7c0auw/Zh5zWB4LAcRBTI0RCpQGaAOx
dJs1klbmLWS3Xd5EYBQPf3LLt6NEzH8I+9PljSxaXmrJGaClwVQPklWFcBiaDNCm
R3WqNF0+saroRcQKsOyUm4AvOqlszt8NCB73HX1ymHY3lxcAWdUkHVGQYlOAHUK1
ekyTSBO/bybJuWiWV+EBGF53uELDv9Ot/gF1N7yPtqMKjQ111wJ4F61PVMNnzmDW
o87Y+REevdznmd+NWx+Bzq2LbROXIKkqErFJuqmZQFJBspf1VIo4n4+r4jvHcdQy
GorbK66OvugU9zu031QzabjYg6IJ14hi3KQA91Xv60Yg5W3Y9B5YK1+YnhsuoaB4
OFOMJRoUScKj8rnCUG7hiFZ6Nv8bn1+oh75ntEu0X2xrrLND6ZBC3yr46TSUFloV
FopHBotg/xZirs1Jah7kbuTfEzNovIhw267cDNBzgLVuSxXiKMuhbrZ644MdKYAY
1Efs38iB+Okx3Un0rKoZvWBvj8xqbTqP/Pw37NBwEEU5L7+ltVNeODQ6rw3VIYp7
CqUeE4z3zKVEcKPeW671gq0QSd+eBQIfzJi6brGQhoOyx+sg4931luQYERorgGNv
ddNrbo/h9Fd5s7El7P+zyHRRDbQJf2JyW2JP0PpdXoJLfIGuLzT6Zc5df+5E12FT
FK1GrAHi1qwKdjK04zqI8rIAkXd5fzQBB7ldOtVOFIjt8nVUVQi2RHTZPZNJbMsa
USpuCUv3GJT7ok+SN3avMKq7vPaqpuwCvLBwivMD0+gBUoufHasP/+UoOrIjCMfc
48kHDior+ahl/xeAwWqjDfnTJw7sr/hfqVQ8lTGczmaRFISHmXt6QhOVWcpkPqcl
V9FAD3EtWNVInUi2uWq5lkgcrO+axjSyFHiIoa5/YvC4YprX7oSgQAhHfaoZ/R/F
w7OdLsDY9FCLKmlljmj8Rs5Bg6k6/to0YxI+CdgUUt8CZr3vPpgNMjKFiPoCorKt
6NAiIgjfy9rS5Ao8/t6NOabAwDsrjFLSSC5PWLO3HGsSdGwZaM3p8nzdRAISKcQ8
VtHiE5O0z5Y5iDsqZiJCkRFIpvkmFCJRSuc2lz3llwd84Bc7Igx3YbQqrdGStm6M
zOVxYgsBKW5O7PB/YPiTcCQNmTn1oR3utP0wt5Zj0dhfYMtl4jKjuFRrR0XXk5Wc
VcejieQWhC5u1s/6+LXXbX9qGTHO4rk9Gr1iitpfUxSsobLv5XquAYaaBIBTR+hw
iiG67IeHYp3s19xv0FCfY8X1ilo+g7W4QC1OnESVv8C4vVpuc1cEk4bwl6iQNivS
y/sUClzS/Ra8ms1flSXkJgDxy3T/H27bklXsyc6ibC+7k6mX0jVb9R7MlR+S4Sy3
ToWUC0c7JKFgCGXfZWhS6uMxxwxmQSif8tn3sHxkJQ1/h9KWcr4i0KSquppuvkjx
PEG6P3eJNJh+IkQogFaKXAAIn85PqvRhZxO8m7yfYoMqrSqdxgClxfhYHPUn5Nfm
6L8GgkepHbC+upnu+JEkf5BtLs0Y3f9d3XdQ3DZKEP/fRYn8mYCmRRJYJfHpKTJb
eFlQ1eXR2cXGHvLHU+SC78nvl6axPrH/dcJXnIvQzcqUijsHs3Lhx644IFRGQ9H9
Z3uc3JEiik2cXRwG6ilwIo5pIBjRt3xALlFVVbwPeU8/k4DXx2/o1oLCd7DsZFHI
hAAjkcO60fO5msTe8Xdd2r/9MZGrxA1J2qkvEVahAepBgQ8R1ES3WG6XeLxuUbJK
J9bXxO/DB+8GjXDUfZCjMgmGYOHod1Vdpyc/VgIfNtep7jOk317JiD2rccb+9i1k
8L8/VSX6u7Vk6H9GYXK2fEkoAtoKx9oq21TichamplQZ73biaQfATeoRCyuU3SMK
Wv9Y0xpPYrBt3W+3xbZeKG0koCCLtx3JhT3A4N2c0yD5GXqID97g/w48GCMgt74q
BTEzObMB3pNJskpv9mye09kjM6dOBbGthPjGGGuY0ZmkFjadRwhQSRa3K1WsUfj7
wLA0+M3sR5hvk2GgJUgFI3tmD+RgfPtkmxeGKE0hII918neucbaRpu6SG+3DIBqx
t5QZRagaFKci6o0whqPObDtrPD1rquVjbXsDMMKvqrsV9QB8FcU3+yjh2LcklsoU
z78ybq3DtOBnZ2fcv1ujIWrgNSY8KsdCwqHXfmz4VFhrxymlwNbRfr+CtB3FvvH2
T1S0nUya1gW4NHyGmHAwLVFSAEjMF8opKoOPlwrKrq42STFaDbgMdXfmLwgrLsiN
tyvDXGsXwMAkQ2+d1iZTfgPSZow3+UgmVfl7wNpNkAuZSveQKm9P0oyBLmCBV1aB
Br/hSZtmNaGGB+N0yZF5LBfoSnZ5/a4wrRQPqzILlvd7VKxuAJE8hZoiC3SJaiqF
bTE+wyxVKDRiJgjmr80M4tlCr19FXym9rQ84Jws3JRRZd9H0SRCbWp1FyQo7juH2
AqVrN4MjAkDViUMttxCwD39XJq2GaZFua6lLsUBcvI8ypRkt1UWSzCGtqmWQJ4UY
5bcWOAB8bswi/yCanPsajV95C79wYMQUB9x/6rria+qVtnbuHOVcqnnGSLv2OmBn
qRS/0jo4LHuaGeXN30fjSPWxZNWj6d7Y+rGmrdqwj3KhF7FIRKwz2LlyfdCqOvsC
1ZHXho53wdXzO2LzItYwWWNEom4IkomD4mJfaIbmtfPIhpsX6VZB8+QnuCehCB7r
fQIYegbhLIVR9sKGy26sZEDAiAi6ZyJC7OvmGqcEitHi+cO8II5pOAyU4QUKodpj
y7k3q7Ejl/+i3flZVcTIuTowPjP2yrn2YqxFxDKWQ7em7FIGNyGGpvisMrehCM4h
PoALz8EMBl7whM75fT6usSwvBCOSSPZZZtzhMJxVc7/GPL/biySL81PG+08UXytW
g+91q4ohqxN3/HLEC2EpfOqguY00VNDAgHpsCZ4wingdoju7cFh8/qlLa0eY8S9e
bleufiN7XroHPI/bp1E3c7JtH7Cw5nz4fDs0EWXgHacd+Ypznx8vUXoSWPcBXBlM
5/tKRxg0AlIEMEVCbG6mzrbsbyb03qmLc55b/TrNUgWm5+KwYbYOrffyCx3JyXZe
ZEt8rhURxuXxjfRwasasWB5nyY7+j2dv4t8l6OIbrlKA0M7FMMVqCOKPAAaoSP4b
cahq6k9nSz69VcIg87edx7Q70MsBC4X2kS04YvcyRjlCn9AWT9H/OGYku6tuweZk
HgjiunL37F7r9+zeOflsV9ucdAYDmE3qX11easJr2YwJf9DO4+LDIOsXOMZr02wV
ouraj3j5utHahmGpH5mR8P1HasGyGs7Qts5S3ERzfnulEjVmKBCyOK8GbAwf2ozP
AFU/tP1IcBrROrtczl/gQ9Tz2K/HnbHeJS/ohbqHRWBKfEMvMqwC6nospakF4xGV
T7E8iVkWRFTyHJDd6ewVYjrHOokgUFm0f+X7SHVw6AsP6pSPBUlNiWswHVWj9Cjp
RPWp69QHNU1LjSLqb51TuAqaxpM1GSC+c/a7acWBEf7M4Mzdo+1PPwgr43/HsRme
fmnIh0mIKowNv4quAgRB22U1/WTFRrILhxrWrLDeWckWP3iHuFa7KdXUWtjmSt2T
Mt0RD/UmcFD+yGmeV6xCjD8G7aKx9qWVs6LS7vnNyT9IxYzgkORQITvzbachm99h
QdjElceG/rGA2IiHmSD/vIrLTBQNnIEXcCBvOKj+apttHnane12IiYQm4JGFlMwc
tW0d7n9c+JOa4W5rVSk/ToyOnRpk7tcgKVGhHT6agmH5ff5OPjZQ10GEtkxiKMD8
JW7bfszSIf6U0iFIuVQe96gXyK84I2D4azHYpMy7u5one9emyzQk42rS2yPtCgqB
+CrUXnjDkROhWP3ZLf/l2gkRG09SzBz2mmZGzDy0D3etFgtVXOjxiQi5EEFK378o
vz+lc7cwWFqeRdSq5dgsXbAgd7RfRuq6wk+BZjjtpIBkhufP/tY6YKwhtjxeKZIo
lveHfndtHhfpEEPbuwwGyuQh5UsRw2wULMhYzLlca91CCit0OZ/iiTzW7aUYH84F
e4QyEvAEgAOdIgVodmBDmmoEv3Q4KIYFLeObqmKihwk9xBUtgsBRBEExjfV7eokV
6gSgBwjHylLNlRiOgSz+eksC8ZMshZgShhKWhPTk9d3JM6jD2Zf2cC9Anlom8AYv
Ad0brwI4WOGUctBSBraytXNkrC5VIYeRNb/l+U8Bp7tcN2fsLwAKSfv4Or+IHWDu
9xlxFV5QUVTIC0D0HKm6nc2ZsSg3xu73A8ZXXF9/hW7xC1bizCiB45rn0cJVT/kW
X580/mPv1cODf2x6xEHixeOxu2sLdb4C1Km7nXYOQUBwNLrgcZepqBmfWMyQyojB
FhZnFjl+6Rlwzham/X8p+beoVjbVfSihYAdA+g1MVdtTsGSO1BZHBLf5AwnNNRRa
qNURb3SLDSvBRiXdB1iarQRQgT74hcgCq8o3vlQ6tQb5sC7VnNL0/nGh17ixYef2
43iROoxrpH0kRcRtZEyfMPjzFsPFiB8wM/umbVruZBwWjxqRNyArInsIbfsOr4OS
63tZ4LV7/xU2T44NrHEgShOlGY8hLl8kcj62JUInN2li30+CPZ9izcYcmQRIYuuW
qmv57NlgVbSKlbJDDzuRHFMsRiQOXegNVCQwmGjNvfze+V97eoqgIv8hG+joeRKK
kdFBqQmHEOr6LANnlNd5sd3Iz8LX/qmXww2K1FZ6z1mwNWw+LeUWvhgYMOjkkItw
jzN9ZDCWbwZR4mKHgVz03PnxP2PN5EcZCGfYXdQgwlOVEgDVvql9Gl5AQoJeWZjq
JYCsawRXVFIb6J0oxqGEgBYDKeHc58ZojptttUKFU/Ak35FNV1c8ayeZz3C6iaca
wZ+9LrexAUH4jY+2okhQa1SW9U17qKH5RtF+RPRp5bEAa6nq3GWiBRrpquyJlr9c
/Z8On5MX+3eu0h96bbHE8tXJgB5dgPFq5A91W4yo52MOCXp4WHozjNAEo4vCCZZE
XExm+0H4FpBwT8aqYNngjrpTJVBRtTrvZpWCut84EkF2twOv0fZ4p4LWLb4GjFoA
vZQjGA+rD0P1eN5n8+rsS9l8rHhufbqPNQt7ouziXEfVVi/LN9ZiMuQBe3bX7BcQ
DKUKTvXmRtWzJkYt2GKWgdJk2WV92fugTBpHtSkiXFWK1A6B4qtmnQE9Kl9RcPlO
bKlJqL04em3T+vMUYKjV661IDOcILg13cjPWtDMvktUDzdhdmbc7xbb6JD4ifoiX
U0iC6GVZgTeevbVNoY43TKQb7sarqDrG+16KMW9qdGgqmpUfitVgy+kUGo1A5Rh7
r/fsTm5dHOEK6POVFviM8Csmsu8VlrcAdFFkv+kI8jnikamK54jwdVV3FwqEscW/
pXvNqlkuXJzvqyvvT9WQlyvZuOUceU3VCRsQDzNC710=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
DFm5/CiL23B7c3uJiSdgA3FFUNa0Euh6a9Ri2oQFLvFvy1bJuPSZ7qriZtEE+iXg
UGevPLh633qutKBmI3ju7Z3l2rXxgo0GENqKkDvCiWDWmSxFsWFQz1BjbS/nrEiC
syVwet0V3YwuWE4oibFTZeTtHuNi2RZGylzgU6Ksitr+vb0WXyBBmRxEEHQ7Nyhn
LxrdKVzJ2Gj6iGUNpculiF1UKVDBervhOe54DKyGixK0BgIPnsXROwb9J+p7+igJ
3H/dJe+sYnQxAwrN4rCBqUxToSpW+R52ocvbWaWBxcOWheUBU8ZtklVoHdsozY3+
uqA3F7SsOakr2iXR/c5cOQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9568 )
`pragma protect data_block
1bliWPzusvlv3VkoDLV9GpOm/NZDTuPaQ2uMF+g///Ze8AAsUJVktA0eKLhyCW81
ra2ERPCVxBnzvaWqtT8uZ3jpLsI22RLLpQtzvy/oe12H9BpRj1dAoHyK12UpmfEQ
YSfinplb8tdf7Ox2PirOQZ53E5ReMPJfrl2kJuDa5yhPiuz3LDXlunDCZlUJHvcH
LK57uCy8LeUZKKhbW9zFbHIz2BUEt8fXsBnRRctpLQbn7aGRrB1Jq8QSOTUYDS9v
lHp5/XbatS5YnP28YUELQ8XFLk7YctTgLDa0fP6RqGmQQY9uz/M7PvVbFV0h9vIS
FvehtvkSjG+uIFqb09GtgMNAR6HoPdJSApeeVkSY7ec0RmbRNHyMs3NZyj3E668S
0r59RSzCikz/Q4UEEnL4GjGWL42OWL+N1s+rGb3ZTU+BasV4hTGMl8z+P9n6RDPL
TWZtMpMHXDJPuH2d7kOdX/cmoo1XmYqnLY2KIw6ma7rig9P3JU25i1OkrEAvb1ud
tCPqLlKxQPX7++nGsjYjNMPKjcMaGwfFWTejUEE2uyGiwecHvlhGPI7UWSWPk2uc
NEp6XAUiLrvh+uodQStI933Pt6Tsne4btmqrh7XOESRFAPq2eCcL1Hjlhq6zCA3e
8daVrzdoTmFSlXeT3HL8Oa2pZhTPBEDME3SK67+to7meWH0KHggFq2dgEWGJo9lv
ZuCKCy+y/4e75ADx58VUQ9cvRnMjqSdggF0hhPx1pWD8IpapV108spKqIL0SZeh+
gmiPVCH25gnrGJYy+wjWJ4/u+YsdUc3xP+ig19RSX5iRROUWobHAobFlkYSOjuOc
Sj28fE+Sk115PLkZ38RoWjNtzP+lsvmbrCmkFbSDBTriqzAJnzv0ddSrSVxTsDab
awmTb02/Rwqie9XX+036aq78g/1sm+EKahrFxkTVxUIT1g2+dNigKwy9mN/6mr4g
2FZTKGfP7AMAtepcdAZZgvOQYJozcFtSZC/mIG7KnLEuJpFohBHkxl0XiOPIX1p+
csMXx1GYY48qvmv8RX9uvhPbsZtlm8WfZqxkQijKqB71joGmXZoYMOQ87/S3N3Kj
0dM3Q3wkAhYoUCSM+v7cTSPvDZITHzAkbQym9AYl+Y06SFxnJOtgdQn1xcS5HSXx
CxjTwGPH+/9Bo/n6282z5VoMhGt6Br7c+Q6Ye482TB2caISmPBIJdPf4JRF53yGx
o+kWkKIKJ53dlLNVAWarESKx5t2bojFyOKepJ1QfSOcIfi1s0eiF8jD+tn08TV5U
VNVO275EWQeVHEqRVaUewpz/vhVdpydi5e0BG8qaxRf3r1pGtsXsF68YrlbEjdwB
onc+Cs6U13YN74DwZjkKSKRXxjZyk198MUrwR5+TgjEjtYsVXJu94Z9thA7QEgnm
GB+kMefO7PSL3GTn2r+M8FbB/i1k8Acb6mUX4jhseoaZpJiiM7K2QP+hFEEZ1mHm
nE8QJPrBMdmolOz1Qz/sgqddZA2Vk+wUCXKlQ9aij1U0X7Jzk7d/LJ7JTq7w3cjc
V09sO647zbOP1UOY0bCRptpYLUq3//qCtKyZiieszFWWcXqw4g5l195TH7NN1t+b
Dxnk5+O8mnMoWUPjvAe9H4+4UzYmT0O5t53u0wIPWW2KCccv9BWJAgk74NZStQt2
2Z7NSWc6OhDZJxNHiHeDEiNAE9IaVkYtnKCtMEweuKaz7oPNAjGh0suhY7XGfsuR
5lBTQCxU974GHb4LXzosaRSyILU0h0iNivobBMa6nYMaMGYV77rijz8WqEKyZ2xm
8ydkwmrmasPEGPzofKMd7b7BocGTmGYo9/Emc9VRENb1bnPjGWDTONaHToMhRSrU
qKjErmlg58yYQKRX5Nkmz+djwSLBa/PzhgJnzc9EWXdzTVIztqb2qHhp9ULmIKE5
6UjCbyKokx+NCdEdnGan9Guq1Ih1OuanvBdqOciIXYjaQlq4plNjUpeXuwt2Na2q
MVzC7XSlzfbc3+KIlfJk4vjJP6Pt77w+MioXx+oIaAkK44NEc5jEnisZ7/eOsw2U
WyDTqL+Mut1NHVLMSPR+OyN9ju4YTwNpzHlH7uO5GQKLbw9SJR9a6rQM///0ncWH
Ttwwc8LrPr4LywWxk+514w9g8gGeM03q8agC/2gO20ASghbdW6elMEawdja0ewol
y789Tzd/glp9uwVrbelIopLeIa6CjPwdL3BsFaVP6LKHulSWxGHT+ZaKxEVkQlXH
nEjcPvciIDctC4n7BF7OvMT7p1WlVmMvcAUMaSMFf79Q/9W5ZOK30vtjz5I1RYFh
mrnUS7xMgE5XduGNxWX8b8HxQWqTWOFJLlKwPk6iGQteD82iaPw9mUZ8EZrZFDoh
SP66dbM1HW7gofFEwyAH0pjamfhS98VLxdlFZGVfzdRPHyczCkxOlLisEBepyIEf
KRWjxo/wyTKvJQQr+081gI8abCd6eks58ofbd1JioeNxIn4mo+7+KWbL2Rnl1dPz
dmFSuWaTQ/5OMlzxHu8JDUTzSzhp5JwyH5mMW1ICD0Dg8cnnSvKCm9Pl+4uDJtxW
lq42B26h9Pwz0GyiNMwFmhzDaNUf1sWUEei/h7qUsD6bYhBqqjuybtDomfJPjvjD
pVv+Ewp4uAey1DtH1xTDYjQhYz5VCxynczoBAzLGbnt0ZC95E9I5ioduBqztTh0X
QbAZZScdq+D9t8RXHLziP2wY3ZN4u8C9EhU0s6m43AclzodzM3q7ML/7VMfE6SHf
IKw9Tw5TRTH3gnolj00XCSF0RRHPfRsV7HlWW7osFvKSbXwd5MmRhgpJB9XRHW4D
5NY2q6ks/56YzctQE9mGPYQRKmLtySqVijqBasxCiNq3Z72TwywmCyz3ef9kmuIZ
LmlAo0D7r2pgV5XF1i+kgWtqEMF7OWsA49DpM8iIJKFC+swCqNXmJE4dE9RsV2Hd
nDnAJZve4QCZdqeZR/GDO2geVJZgVnblupJSEEC9P/+HqffKjHWZM7SALPMu1Zzq
w4ypUwzCRFj7en1CzNZQZqfNewBlpgAsXPt7wpq2KoFwYgAGinkA++W9+bVVg456
J02tBvKlcRrrCobOgLpQDMyJiRaPNWKUW2cmcWjbIbDs10RAGVmschIrJBqSRgDT
xtYDTVx7svDXU/L0N61UdCaRrZl7nzuXPG1NIEjvCgK3zhIXyQy7yhD1zYhQ33Fc
6oFGQBW3Rs3r0yTKfE7m0QE9kAKuRnN9Yv9IVhC2IZ9UmANmAEiYzvGRHSlM/rLD
6z88NjqiXkdueyl7ntkSCF+asv43Qy76ye3tGe8EqXULtDaokPuTqlzaQJfSkv/W
jAEMrhjsrhu6RejWTJgx6GyLh8quHLFpqPaF/nfnn7lQI5l9XRAsKGIfFHqZ8XLH
+G9whOs8EIWDs2BnJsgal0Mh6sCMavwYXn0m5Ao2/f8DHUniKyIAjG8dR8h73DAR
QNOK95TrBZ5X7WQa4Vt4JyzNAuqhT+U04cy+f8/8A5fBxnDOqCrGHYxEFERUmD+M
oFiwxTmsNnU4ohut6rJYYb66PmF7v2cmEGhHqcUuWJEZfV/yBk+ykeyTZOtDbFXV
hHhYuprMD/DCJtGi5wQp4gcuiOLN7cyeF3vEYj9q90nmXnhOedx4zBLC0Pc1WvyA
eU868dg2+W/GUPml9Bjg52EdXa3R80b6EiKzlof/bgt0pXUKwLic1hHOhV0N1KgB
EmU/hVok98SY2KCO8UoVKfmpOiDfgtJkd/kmDL7WIPPvnjM225qQiAk+fP5JCDSc
YiROjrHy/3UJYmXe7QDfGKWf+BJimAMqpMkERxr32mIeuTZcuJ/1bQlDD3ixekNy
fxzi8dlJB2aPvCH9+803RuSTh0Zvt4nIqZEZEeIJg+urkeOPcF2Qrb95nLxW7FU2
FSSk7GbIsNOMJ9kBbK6xSe+xE8BtJoM6HKzNRmh414MRnuXdIr2ZWAH5x8vu8Wa6
1DX5VTTekzZUbYtygMS0pltZH4xN9Pk4XEr27OaKokxwidXVl6wMyGRDZyWtW9OB
RpfpdnjemQ/V/p2aUfM3qDjawpBFQ36Sj+c0Ib2Ygkz/3OLvzV4XnfhlKqbi3IxC
l3HYoCDczo9oEEXyvjmuJxoCihVfEDwZIqkFehs/xiRBBam93s8ejy9Rvdkymiwh
jm/v6y8aYjsVqLExrHS+uydEOPzshPx+sKPNPiDYshZT5eqmZc2SRhJDUPCUCJnl
6lcY8Lz6usMJECX8SywBJ+KLoueEMCsxGbR5e1JMwcAyuNOmqFAVbMJcwVFCouyy
IZLrHIrzT746eTfTv/gHs0KqXz4sijVmBNR41TS+cgxVt+junO6ixxWFcAx17Rn+
Q/7/LXC08mmbgJEoQbsRDf/0Cb41ONej032jxiNLE8Wty1ZsAmOmfj7bx+/+QWoZ
OhZ/wWSVfhQhGxyeQpmu2Mxvp7hY0Tdo/68MDevw+zxUA5ULAKnPwQvMjOget1yU
mZQNYMM8ob8O+Ne+AfdtTX/3DhoZxw9J4THmaeRN/EoshS5MkUPVqOS1qw8n1iDS
zTUT53GShnYAsj7PO51CtJyYGwiSIozP5A0kpFnLuGGRaco2IFB0/NsyJSngwrti
3vFtqjQouN5X55wI0Uq9WOX52P1dpIeoKOBe7MRMVRHrjLSt1z+Qs+TJShbF2CdA
eY0xPIw2JPrT5N72UFPmRiYx5VU8EZp9Y4SgKA1A5QWYXlxcQvZgpe03239hGvTZ
ZU4xsobtRTi7Ubm+pCvIoCuLIvsmlsjPvVKGfsuiNnfy2RxQb0fjMRsabBt3SriW
a23zcCFRqGKzUXWerkzUN0gdlBUhTrx28hSx0u/xg6Ta1xnHiNLrl6lnb3KppnEr
sX/rja4it076Mx1GFwkuYCblepSBT+T3PEpI71zSwULRd3G6pV6BZHWmXD4fjXd2
qNQZszslHS/glOPBsYRL+2drHkcsJ2xG7GN+VWPG3O2/UzI1aB4GMc6WRw7VvqUl
d44Fmy6rSRFSvgmwuzKqELv/SifwRlYFphfHOnKGXMXvEtgYB5rQ/CRVNp8Q0BUL
yBCA+0PO92Pk/hv6sZ1povZNbEkruhcgZP5vgZNUVAcqcLmAKadk2xarCBCeNExn
ntHh3Hdvt/Vr4j2soNZxzqdNYhlSN/tzWyprSt+fGXhOISia5I2zU9wVH3xR9cCy
/35o++1LUPMfM+DrcYByXX75aiy/hWAtStrBs0coJynhxqtTjAgIIVNQNHVmBSQl
pvAOwKzuw4HqyqQ4tF57rXYtdT063I7/5VSM5wNgqho299C+FhYKI4u8fXYdje52
BwsqrnsgPO14UB8t2dIiz8/Csc8KZkE2aaD1vZwsEmIFv8J2BWlxNhJPpAvWkiTp
q+hdN2cExS4/kgZ4wqxbdNig8c2+JT/4zusZfc2UzGdiyUVzdH8iGgykI3nIjQev
M2593GHlFgtOYOwlFgvrd/YcKOVUw+vW4otkg8fVkCEIGcs0lSN7pRaXaEIazYsY
IzA4v6DiNy1+d2S1oHbsQlPCzaFihZzX5fU1Bhc5iIZ9EOQXy1iF/WvpJHcy6zAo
2824tIzPhDZ5+OSf1PihcXk5nl2h7eUXDA6lyhioXb4bjb1R0O9g7olY7GJfkS9k
foAT17P26mSiVT+q1vDJQOiuCu5lLWE7tE/QlYD4Ywb50P57hl+9NbSaVORY1AAG
OqjnprcWQSkIDA3vo8g+u0XyNMYR4nrl/94CHr95o7q2QHYMl0yUErxy6AqWTPPZ
Gc5V/eyPS5HTQkvpyE6Nr8nNkynrADiNSlz0QrbnR/kk17tg7cpjJVwCqkJX4mDF
i31VKD+LpY1SUzBhUp+2NBhj20Mze7WiPIGRC9h5d2J3taUTcH0xO/+c9S73ttal
KIKDF1sXiySye8m5zhfZ0k/V5fesn9oUsPUYOnhW7E39RvuiRzxRFNuSNmmnjwOA
06dnkUHpM+RFDrkpFbZayyakCSQtHV2CIejigRv1YbRPTGvzbxZBzadbVieNTkLj
6PtaSTw6Q6+uX7FMM2Xic2l8GtUMH/NjbI82bheP74vgQtKyK9cCjzGbjLGy4n9p
E4628bGSbL30DovR6LaOab2f6rqGUK1pBkOPERssvkTHGVlkwFAtHgTmcvRxMcl0
oJlhebNYXo0ieKrhS4pFhrPFaQCZ7tiNFaL9trkeyG+DmTPzEn5YlmSjbiZ0HhMr
7xoI3850mx2BYvsGUexHxOO0JtqdMfttLi6zwuenZboxflBwGPRQ5rkIhhTua62k
u6X0DoS+YsQOUgD1Uu7i8/1kmd+Dwp79ZG/lkfUbymgv3SZCeAQI92lasrE0nAfz
CgOFZ/s/ixenijhvkTmdxxxtTBZdjJrU730Sk6LBpuSBwu1us3ROGOW3JI4nawhU
Iu4bU3c2GzZ9yhhSSDgYJRmf2YiBo9mwyPwkxW2OpWR4eFgBc/ndutDAk8jy+U95
WRJq49lr9JkKvCn7je8Zsvpee+M0YanzgnVpX7pw1pdTo/6ObfDpl21HvfSFb4P4
YQjGvW4/zgpWk3Za14FcPi1YFvMWob0njECS+pqUuMNKI7Y4yk6vrIha/HHKQXTn
tzinInGFbuPG8IVlf/bzvRR0VLSNj/rY1VajfTtgs7d1ydUCtJreMsgVd3bX4PT6
DZngAn849QC6L9o4fdItX9FpV6WyAaSSp69Qo+KFfnujiR+I+tDZevYSfgp/k4z+
fhQ6ExEa8OYhlTS8OYP3wSurqehjq2EgBxpKH4Vr2F2eIGFv3PKRiZkoY3eH7AvQ
bYcMZTSmiSn5i7StUd5eA2M2hlKdSA1hEn4mZXLsY1E6LXgfts733KbxN9N4Wucq
snyiHN1ODWqm3Vch/ESNud0H8TOqiz3tuUZ1b6vNQffMHE8CuiQVkzV6vLLsLalx
bQbChgT3bcDKv1oWP8HnifBZ/aHdFay7qNBtFJHG7iZoV/n8+iRWYCQUhnDyq8QP
/yFn7XJ8SQSwwrxcwzi+/Cr+834Pj4i52NsOtwyjIrP9xWVDAEyXPG0XNSZfDR3C
q1DDrRdXC7foCPvLRHpet5W0L0BUmoSuRh5gp/VDbRe9wNyp3LldFitNV5RmuH5e
3PYXU2WH/mZ9Icf+mXCva3xm52ILRrr5jvpDxMgm33joJSCpXQ+FYJbXnOr+AiNI
4szvrtXpiFS/M+0SuZTCi4RF4U7o9lieRv355NwMLONTJYV6Mainahlm8JUhTpnS
x34i9wgFx9xhm+ixPwzWBSZu/P0RJrKNpEHaAGFt22CBuummErL9xZY+feUmdr0g
fReGzzWkzoMRh/xBB3oItz2oMp8JcvjdVBd5EMqap8BWCMyDTxEnkch5/yFvrJw8
vdAPMxjFLKCiDC3bde8mZ/OPgEwdU+5hKsBFDtD4n0CAuNfBBymn1FnEwclE5xz7
PleYU8JOTrKJq1XeYp4ME8W8NYijCQjcuR3t0uOAUynRVPhItZtp8BQDXuuRiCTs
UzJFqECOEvhpoYbHdBG7m/BZKUxUbdPvIbAYNbKt2lb9bn5RKjCGhNg9mKRJNYBk
qLEouMltLv/+3882AiZtGaoVS1jKv3vfMjvKMjkTGxVyAioggidDVlSwH0RSJlj+
JqgsrMK1rKJPxha90mLQC8Wgr8txCV1N1S1epWqcmFQzB2lQUt/i/aFXNxKXkDIG
csrfnoaMSXyuH0KENvfYQC9hB1FMhGgrUc4Cnhagr29rcwGS1PwjphSaHUXDyl5W
rz8hTzHYf7JKTWGuDaojA0n0zBz6sDshiPLpHJL8GWUkZzg7qiRf6/tqgPVomKIX
5+rWrlEojcPPCZydAvAfLsDTjmnsD+84pHuLqXqnZiAqVH1JaU3OZFjBU+2M7opC
UWTgoD6frzgCFFG9pK2E9P5MUn5Yn0+f6JflJKn40/5Gr7XU3f0H8WqkcEIrsW/q
FLm2hxB6icRYUhm97mE9spEdVGxPyks/4rUjgIp4JXssnjQR6e7hBQH2BR2ms1B5
kdiMhVJeCrlyIjIqTbEaI5ReqRo8P61RRrEM1MhmFiqmVn0fwJuNZ3OITq/lS4T6
kBqsdvKSq0FeAG0pYR38xuZQVf4mkLnwdGeaVGuzAMkBFoaf2uKkghsX5NTReAgE
B9sJ+a5yH1gywlll9V2xV8Z/eeVkd5wmuJvBxoqc7JnnJjW03AJSuda17wrOUlci
RweGcdUrUmPdUYLl2XPJWJkC8JqHIESr0Dh/l7kue0gIqvNmRhZ5cRfiSocP57wy
TLMLLDH09WozxATHhJd/WtKMdU50E02QMx/P9+EA/zALhkkxW0sthBBJn6n/ya3M
JxxVxs93vELLKzu9lYIuXs6j/N/UJ8jiP382JG5jGzMuDXFCH84x3XKiXk7kih8e
Qbwn65xDeYOVTliv8ZFMLnirQz1gB9Bxuoeo6/l2MTeq7Zdx6wad1kxGA9TEpD+3
3+E41efawp5Fx4thhyTvCEIiVUOtfaI45ghD+ypqVT/Cm8aWrE46oqnBuF/6URc0
rdqiKvOXZo4t0uHqTPmAyuVfLOoHdZZSeiXK4BJT0dzzAwpOuJsxQr2TOvpQy2L8
wCXtdorFnpsqx1IHTTVUAQs8ODRPxSI6g/cJDvaTt7H5PhvyCi8rfaZkYOfB4CGK
mOXjPQl48C+2GPt86NJU2Y08EvUtlqEbBJJrNdLO5c8/0p3be7pYKAKwOuwvN2eI
eKVwy/lhdzD1JY8UYViViMEF10ErFN1EG1evvXi/AGzwO3gslojc5m81oWOXSaYk
miQk33X8eVI8hORlUV3ud/ha99diqGQ0WQFPiMNY9aoT29PE5jg08RzBMUXy+nZW
CyPt3cuuacmk+VNvKpcLP3jpssguOUtynNHmevlMY/2iXasyGahjsOj72hrzNQAe
3vl1+dXw3ADyxDq9Cp58dvC4SLHgYbREQ7tE9VjTaGsAwx7zaiZlv6E8BAdR/X2x
uwx1ecTB+7YQx2Q6s+RmrryBSYkxmlM4Hi/03QlNdfJ5CJISOCtakaKK4S1gIMWD
2yYb7rP5Ngo2Luk/xzYVydgYyztuMEhGzSxxExgxz5EHuQuGnUGu/IpS08iV9DRD
CqGcSqwWAsNc5staNacylxi40cUnIt0oMYpc1Q4R5B72NUl2kXzxUtyB+O+3GuMU
8BJdrQx2aIbe38T1g9/Uavoa5VwioA5g2+UBgUFCBBPBkcP25mt/cF9daDYP3KP1
wGRhHidkFZRVqcnNVYv0ULAIWFKqVRGgIPZvjdOVydHZ4zcgAc/J9vfC+1XWCHtQ
8G82ifNgo5CaIJN3OQMdMVvjgjLiQdnM6g3sd9QzD38IYAPgGgtSWTKheCIl/96R
5j0vkONQaeWnmxoDWbpEg/kbP1nzvVhgkipZtUjLvxAwumrLq+5Yd+lIHXlTM+i4
8JSG031PwDTQU3PGkH0ZBSzBqMXofygJa98mT1BcKMB8duSOvB7Z9p/Ymsw5CG7d
9tl9lDSCzjc1aHK/KF4BnFzwOJ87O2EbUbXcfET4p68jbq3SpNC15a+yAlE1IiO7
2y7J21P6xVSjIPn6G9BlZa43x2XN446zLZGL3pDihGY8jEXng7/BbhH1mzcCjDtJ
qzLR5hVBfHAermgH8fNHn5d1hHmqc+HzV6/6u79NavEkX48BpYAAr9NHSMdWhVtA
72IBRgyg9RBRYwM/wJWFjSNvS8PGEFEDGjUM03nV43pvl3T3vp7AV18L4iukQLNH
/DrhUmNVq+eHdoNPaA8/qkbzCXzVlRmAAeX7GF/E3ydLcB5rGqrR3QREBfWYmVN4
wUDlaqNUbfYySHc2BSpWVgE7gsvERlIasvFwiXWhDAe/8MW6qpi14xtAXIVPAfDV
O6XI7sQA2QBNQNuv47KcdjzdYmdWC++XUpV3Na5xfgr+n77XySrt/ad4mtIkgQck
cNX0JGjFtey1A8V2i+J8v4L0kpVSAjP4DWR/NWOlBnIGcY2naa8FxHY8miF+uY6B
8mx2Os6aO6/1UvDyfsEnrHtDQcGYW/j8KGd8i6NtwW7eRCHmPxA2/XOZe6kAwc+Y
UqiCz31KxceBe1C+frvCBSX33Zc4eAQsNiGER8vpSdW/X3ovqGZNFg+cFtNe10mD
SQ4kVscq9WaSZW83jFkk33Y2wgpBINYXsuCVYM0Eb0dcabFIZsJPn632u3Jlc4td
Ww32l50cvXGitNEeAb2zIAtO6DW4DY3W4IfrpJhvEa+0+EOkzM12qTuiOz2Nt+zi
jd42UF36H1XLs/TI0jDqwZl+9t23ByQeqNMDvHeFy8tFHe/69mJeqZ55jJqcArSg
fL6RufiPVCV2mUuNpAO0fOoSjFc5+KS1LdavXVVHsuhW103aliCx6C3TvLTGUnQx
2SniKyQE6GJ7qUsa5lBJ+H8GAlOSa/tgH02JWJg/adpn1+dXLaFQzCcbHCHNuBIS
mf3xABO2UYogcU6WBYzAiacH3aFbX9S+UqxHHXCW9yUiajwUzmpjQ6wzwntjjr+P
vUTgZ7go32zor2NclBev0sg3OhSLddyU1r5JXK0aYTyjpMKnX4ep+nNB451hoDLX
0oVBdNOm06DcfrRuy43Gy4BVFZELpfZP+zHfbsfR7H7guMvX6G/MVzwEyl9+PsHM
hDmGQDX+R9uVOYzBnQWZf8Bev23qcM1JlZ3DPzRB5SqqFYPa+appoNm7ICk+JIIJ
46DZk4V8vqccQvivDpQ67Z9M6OVCFlnLd7wDlyd3jI0dBq/47v7tb1cef8/Q2GrY
EHlIuWNAktQIssNGtmZZXzQuVp2Y8YP5M7b43+7Tdv0vdOGE9kw5+EforAQ2chHb
mJTFYHUlKNs6W4g6w1Cg16EOBKsVGHkYeY5/l8W2lLzwhk9Xj5HL17rhMJ1x1IRd
K3lfZ2zWZF7mFEaLHpdj8SnTnNWFf8nkaC6oM5NPjcXcve2rjQnZo36JlEjxdtT7
khorZRvTaaZbMb3N5TlX7MT3VXCijjWOwJp7XtXWNw1CLc8WTJMQg0AO74KdESEo
NtgU2q0nHz0bfhikrJbxfmZPqxt5Fg20kkURKtlLjvAj/e8WoGJSLfVj7er4ZKgm
zWLVBvXsjRuXib0PNt0aWIzDb3NJGO4CMmcFPBUsFZ5LvK7HsUliEuXWA9CV6DxO
+QU9D+x7AUhBRsWifSslJG3RIFseG5dKzW7K0Em3RJ/FiXEVOMF3ztdTENWa51oT
luw4yy6TSiIAsms91uxJdP+cWPJazRDiX0Q2qsOE++hOJhjYS2EJ6ulACgvfbXLn
afc6dxnfRHiJiNPvx6z7C7iFJgnhLI6yChqN8+J5GWNpkiI/OW/OF75+8rGP5E+k
/X1UahuaoQ/HPMK3Kjzs/GmBD3Zi+jQt4Lg8TbRJ1wEHIv3gNbuTVQ6PWjXZy7bp
urNUtDSN5l2YFkhzD75uZbmH3wSDvut4gDFixZ/hWom6fi9ejOVvHlv0vzMrJs8W
/BXFFi8qA9PL7opzslabou31aUwWvq2a6S+OtiCL8upp2gvhaTzU31Sooah2HVxx
uur4EBEHp3CSPNG0HklJot4tlz3stLStv1MY3N9LwU4XMqOPkXR3BgX7Q629WnqW
RoexHh0VhNpyMp2DLMgpEJklEGN0oHlTxf/aBm4BA3XDoIQXDLaBhtIvjF4L4bix
xam7SMmCcWkd2lcNRUGXlUgpJFt38G4rLZSB7gbwlZCawZ3v7b+6tQup/y/u4C9s
9NWpyg+AvjXC9yu0tGojCMeXJoCffYH2LHPZrfbt13gjP8uhrj3/PB1QtTgr18A+
JMiJ49+/drv28jaIGmM9SeT5QdONlbUK6jzy1xKb+TmXhNBavif7DH2zTvteAukZ
CG2x2m3oN/lEnsX4QTc52GmT+Q61n8PG/2nhjqlS9QFt3CHZlCTIMwoHdO6uf9cs
9CRrKmYO6aMe2JEhdMp2E9h4laZQ6ceJAnnr+mjeEZIwk+lg/MB/0vq1u5mxNbZo
d+h6YjquDAwH/BcFP7rC8+OqcKRwH++CVg8psy57byZx/sys1D3nhVftKs/DTn6u
DVmeir8Mhnrc5fzmkcMOFgy3YpJNhfjwbFxm0TXISpbV5fNj3GmjLsNnRut/e3rY
GrNcKD+aUGMYswPsCRyGbyVKH5DABGldYLSSqtIZu8wsv4/2lGyM1XWo1WQdymK9
7p/VqU/olxLY3AnstN9m96dNIVVFxrCXig1eQxCZhS22PlLge6evmp3MH6MBEFfn
Xpx7nYDoYGhdxLHOkmx7RR2oIRAPp4Deij3kk7UUC/qh4An29PcHrFOf6PMIUfoN
cZPsz0ySEsUavgwkGMPZx+2pPq3E/YNcgxlC3KpeVpqUYTWGtU1xhHC4PA2Iu6L0
sdj4zhe+rr/K8qkBiAImwGDvSi9Pb/N/aLbdPlwhtv0OruR/SOakRRu/C0tTmuOI
Hnk7ThIsHHlMM2VTnI7VDtWLOhAty7wuKXTRs+LLvr7ee/OuYrdp4gBZrxYn30nl
5taz8t553NGgeAUHdRu0LwIKXwZHpQ3LgBTcfKvF5gspOIm656bRg5ZVZwlDQKte
2G7vESJX6TL2SFw/6J2TnI/LZ+MQR15S6gqcKvRt/PdvMxkgUsmaCG1OEdTFzxU8
xdcFdb8CA2Hw4yQz8O6vo+t8+FqUYcLMXPJBDu3mjw4gq0+X2k1wUk50q5g4HegV
i6yt/XlsmrbF7QDnuNVNH0/QcFrrPEKra35gnaN0hBBw6v8XIhQ6NlUTpKYCaH5D
B8s0HrEIRTzKvIoeTsGfdA==
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
Gw2lWPvrEjGtglXDFE+q9BAhTtWDw3abB9eBtp42MCM3pvNKTYZHlf/nQLubAG7N
VHvZcUIM7OXAbEV7lsglBjw6SvQF5150RnWnCArQI03q1AHWaLVO7YS561GA50l4
PXRrRBcY3KwHAJFM+g3SWRT6nJQs3eaIczhFbHaqGumT21KMV7+oqscUkbsNia0r
SALcLLd0f28erslS4oQ2Px9Kxgx+FUwKknoLrYHqK0zYWCr1bJ1c5LbV4D1rNZka
DHypyctxgECgwboNA6Dqeie76GZFZhZKmRpUz1D8l7xSR1MpH1+44jinbwE2AKYJ
q7Pcd5iRArFDmVQudKErtw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 3440 )
`pragma protect data_block
T9jIy/4b7kmCDxk+x+unB3/1tEOE82G/Xu23UC7+2ClifesM+ctFujAa92ujSdnA
efCjPrkB2b0K9Kv/hcY/uU+1qMd3s+6GDS4ZSSZTyZfLfpSw+y9MXhSYOcs58nxa
0D9hvW7QdiGKePxor2nNGPIpQ1Pz2C6wALgILzdhc5I1VRx30CFrt3/kwsF7m7qj
E3PNCt4Khu6amCAWq9iHs5e4LH717OZf7CUrWf6X1w/A2+ToTztZLqtPmWhSOHJ3
ZZRPXTVlOpt37dquxHqm1Zx+EgQhz5RSB8dtjFrItUwKNq3haNxRB7+rFAgJyGSl
UlLu7nmayW4v35NXH/DwDi8rI9mPHyfk4g9YJm1cecP3d22rt1bWirzp0SruyqUh
VG2It8f/F+fArH8kCDDRrN5lFq4SucEvNE7kbGievMhRqCCJWCviwBW5asqCqC+k
iNL5N7l4Z1xpSBkW+gdI35Fp/cDMrVdF0zG7ftLFMuIQQiclgqDI5EZkLJiRULHC
k6zUBQWWB3hh6byzMci3OerVr2m55ZJJIsWaooOcOmvxDWoZ5BTMefslamPbmDFl
0458PxpkRMTghN2fQ1wzhnM7c0NXFxwadlaPH0VX7HUc2XZrr0BD2QTBN7RWBmRY
HOwodM7LBnA9YgsId2kuQh+p1QYSmaGObcBWAqAU9zlHxM426gSMrTJgf0sWGwyk
MlGkApLIIBYL1iFy0dYHR2YeJTJztZubw2848O2H7Y9WHolv3v2Yo9O1cawUREjZ
8JjmkFKxO0T47Pg9WuKTWThJpXWwk29SxenBFYYh96NSENjZyaQ6zS0Pb/OAeiFB
I11nUGPXolV4Zcrm2lEeQG69C0Q7rlRrOw/cXCfukHF7moC9SmAsGsHA3VVOCcpt
AV/lOQW+sDX1rvrelFs5TUliNdC32jEgc5/htN34EV+ovDGirx9RuHn8uTJZijDM
iSt6WInpD0N3B5Y+asN6ek4L9g5uhWo5nZqBx0zOWAwnQ0KcsM4JTSYaoHV4ylH1
zHKV4oD5i9vaENYHbaaToEnrs89QsJf3PpOim65uu0dzYm/GQgN1RsEHtkqUL2mb
X3OwJ5gwVnxCzg530U2gTqjNMlaGddBq2oeTRO+VGyu8r2lZFlb4xaJIhfVtemWH
7Bcg453vipa1DWKTT+NkYwD9diz36jx9fWaru+VAUEl0Ng+uXsh+sluaMXHmR8yQ
TUd/7LA0mRLvabf8Ru44D9UbUSaq6CUYRAkHWPOZ4cYF/hDTdESPZz5dZ15LRRO5
YmKN1O79A+K4V5Ko3JqkF9lVZAauRDG83Rs3DbWKRXSc3azjmmXJAsvheOFITt17
CXlrHSbZKbjfVbKbZYQEwylIP+Qoht32ECZ0+SSJFkhKLMwZhZcohWaIR6VKtTWh
KfqDLSCa2cXQQ8pOtaZZqrBRTzrwHzeuEzJyevZtTMv/mneA6lpO9hlG7bEtk0C7
7p/e1oCuqEwcyhGs5Jl5Xp3oRPkC2sq7YoVOr8tMt7zVK+5d+e7xLqUr0x9cl+Bq
6rsG7jNmvmcOpLdYJaAnc6HmydCNKSNMscLrumf+u/sOY0xZo513qIut8adYg/e8
HGqsb/muO21lhVuGE0bxrnXSqS/Pb2v6WZ6qewAZW5uwg/A82VEimnw9cShs27LO
+sW2czJxibLb1aSYqyQ9yyrBxEqkZ7mo+bcR2LY+ZPyDfwl7BZCZvM1NViQhWrVX
l/8jQ6vcwSYvEiMajvuUgRygnN8/E7EnkjCZ/HLA/miqajA7ynMCJifovyFzKRs9
wcRvr4JiDs2H4ldj39RI//p7KifIb1EyxOp5xr1F9jYqXnw+KWzgby9lS2xL/Oj4
QgRgRfPGp/xB62j1vYKGtxZiJ5FejCdv+/up+ioNRDo68A5kfkTX0QEPxCZl3EXw
Ds7Nga5XnO3V6GajmHY3BFU/HFMZsSGSGRbLujw3R7cfFkJ4x/uPXyNjeumu/qMp
z5+faaZFy6i6xFgJxglZ6NYebol4vVOul480EoIfVLJmGY8y+0W1oGBrHCy8H/tA
j6UKA6R0tjdhy4aH2E/qKXD/C9A2J+n8SMbp7NOkTzOqXDHW0NTDutRhOx9jUbD0
Ev9s1r9Eg+ij2I5aDF4oEuBSr7f29EeXO/HgFNNn9scDVwU6ZNBzMoj3qLdRKIXp
hYf/hAIwJHp6p2d07fLMmGCRW7nKvOmdLV49ecpw0O4XZ0Ua4J5xpO1W6BirvJOX
OD8nj1ap3rAY3PLmPmUZIbx41R58/eG8WmxTP24aW971UZ8nXBeh7I3f1WWR2iYT
XxXuzNc8XaB1dDYDMi7EskF+H0D7lizhrAgAuBlcMXRP8cO1CMKEu5KEowslhaQe
LNnVrmeMFDebjoDcD26GxujUOIjQS5FCozuZAJJqnCU6cqQWTz6727ljI0PJDKub
XfIvxU0TeHlZUwKusGAUs2f75y4HmJybupd0lnAnMT5vCC3dQbXRrEKeRyJ6s7rO
G6ea2OB05VuOoYU6DkJ2ndZFu3pkKw3/kee6+HV5T4GhmYmj6yhUKDyNIJ3w41bY
4EG93w1V5GDwFR8qqzf2kHDVmYLFrRPbgl5WKXXlk1dgOfsUS5eg5Koq+MXp/rd4
aFWRDE+VVdkFqLkCJ266HYgYM8330dhS/14yFJ7tHEyQDn42u2CIJ/cnOMOucKnc
NowRW9jhHkzPWfVtZMrNnNMZ8zyC76e+sCxix5PnKj9wsHlw5FaxGcdnDfcwuBN8
32Iq7d+BtDnz3KPpoPq9bGGZh6mo40ZLsazUwpA7cnT0xdCqXGiuWGqNVRPYDnPp
RyRDWU6kxQTG6uqtA8G8MVsi3cY/SDPBL5dYNpFsGx+OukRpuReUExApfP7xuBcZ
oCfcaaeZ9MD/j/xNQywcjWdwdMlJpENefkiTrPrK6tWBAhCA/B6QHDEP/S9sRyZ+
euWAsQAUpkyyndOxPiWLNHENMHYasIfCYYpwIloFdWJ3E2+VIq9xrDeQJ1kfkm4h
L/rtTk9cygLn8Cq8b7T58Mcbz1JorWADT1CcaJSGDsTF4uek4TvXyPkzfcRJg+Nw
5rhQjPSqydlOSA1lddDongOIErLBkehe2xkMFYZVmRq3yzIHrcUOhIUVMU6bPetv
Osg4xNrN8XClBna2Y7U1zm7+Gd8vRIqn53nsUFOJNIeFi1zFRcJjvIzsjkYRh9zC
8H85wJ2vqFf1E4Npa1JgCoZMbeeZLNIqfCp0KnsmEftOK8UqIZrXyttO0JuaewcA
K10f5T4eVPjCAQSdGYE+rKYPybesLpJ6d9ogGDzTfw+0QNby3AgKAFBbkSCowTaW
Bd/Qwkfy4oKNG0JcZhJZ43y+fCeMY7mWZCs+rhdoopH6b+PPBuWVrducyCh5jcJr
mw/1AHfezyV6vXkvSlMPS0MoxbDSKkXN1AjOpEt+stbQzNNnMX3NWVJCXDwCXq1O
ACMWrAdFyL9meKVyqz/8RME2C+8JGdAJi5R1bmQhs72RjAVlz/TP09P/XKEDdWDM
PBVaUr0Oz18Rpy4ziZwoMjfe1313x+WNsjcEpHUDgg2sr7Qf0f8I2/kVu2NMrvhW
1KVJMgmqEivkM5QZ7CKQ8smqybdPk0lQduqtvc/aIzKzgh9az+rsRYLcmB2C7P+e
a4UgYiU0ssiCxKX2rDCchlYsRAmS+7Xg0IDw69m9M2Tn8qBUrT86WpqIiEBixe/8
IIsFx3+W75FKd2r5QTfL8UtpEfDNmWmEsMOGf87OD9iDU/oGNtmraXgCUtWhfmAT
4D/KihD3Mqk1gtB5yTgfL063LrTLzjgqM3TQ3Mu4DC7iFBf9hPNjT7gYi/cZrXB5
vJdlxbkDABenLa0xLSHk1Uj8tPE/2+w63DUkZfNCbacaEfrRfloLqnju/aeCeReQ
0cZuaNwXaFITj8Y9PsCZnwjFHxgGDvgsj93mOjud+FK8iGem1YR3keyMo76/KZuJ
OYaW97NjK4r44h0gT6unzRXr+by01KCYBRiDp0QkGTqPEu8DxD1dSCkKUCj2T1fN
7eY1Y0dG6y8yUtaG238OpN6Z4kqN1pohcyk7+gs33IV055p3b/ITjHLD2Q0IS4fv
gnKbeSzfFvhh/zPmZvZDC5yx5KGS2psKs1J+Y6dQKI/8ggVwOQA2YUzKUHecXtwu
YmRlMLjhSeTvfGFw43pqv+BtfsgaBks/J4tUJqEwZHRm9GHqeBfLuUdlRWCO9Pe4
TfhE/T64vvj2zrlYcZmt2xY/9iIEEPXcyXbxhRVM++GljX7S6CkkjYvi54fjhcKB
ijnvDt7t0SrBJJKbR2j/FxZcvPE7GiHPQC52x9JEsGrZg/Hhrge4PEhoaDjSFzcR
FrmF4D5kjNLQKhPoB79KFqkyDee0AskHfm7wBFguOeH5xaRAqP7v8/YsE0tzPHbj
foAnXzKGbkXmwyBvuwiVEHbDxKrZWXtfwSgadUV4APncWh/O2IooZrax4jNW7JfM
+00eIu1fz4ZjGkGFsaR/PdQE55mBNmia/c9WO5vKeQI+g3iXlVQ3Vs/oOMZHl2ez
m1qSFpFFXpUpKO+8p3aOEJbj4grt9kL3WqRIpG+INxo=
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ns
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
HdF/57UmhEj+kkIKvBjv+za6Afz/VrtcacrnZsGP3Vnn+NXvhTl2Qa/Rv4uhV/oU
z0lDQ4E5JEg3WBK93QgstaDRxLKdhWvV3ZKsXl/GM+WZTKzGGuTDFTNS3U107Z6k
EyQrZer6yqzT4FJVMC0NL6IvJpvFwYda+7gjH23FyYf7bwFSuAdISSiIQxqq2qyP
yAWghflDYv1QnEtcpIn0cHFks0cEuQbrDsyEGVP4Ok+hgnrE7zbIpCAks+c//ryc
VwxQ3netCi+apmftQF95XMHfneoRCDNHEFDTrCGUzTPhgb/SzL8TS7CzpiOIMvJG
frl3zKHvRfQj0T/lid16Xw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 27072 )
`pragma protect data_block
b0PtgS6GJqSGFi2OquCZ4LH6X/d4YgFbMwlfQI3sPJeNQJANYICBRDuP3B/wd8Wb
C07cemGJPuu0wOzTvRG3lF8iK6Fxf2AZ0DrP1dxR9qO7bpVOH65Nrr29sAvO5YZ9
Pn5lRDhzI18hMnZrOKHPXoJ6kKYhnX4S+NXTXb3xjEheGsj+TmOJ3fEGkVl6Ui8t
Ght+7IY91pBg61x0vm7IywUWKfY5rdSu1HwhELIPWm2yLXlmWAgoN4Umba+M4yIN
9MIo+TtzwbpS8R0dTF5+DAR1rytb4G8xszKcZi8ptjpF/qTypJ0Gz7UJD2bKLlRS
56sdmIFXDLh1/NO6rjfYUTMLpOGdV5ezRhIJgvPo55pDzsw8Byc/uOrLS3tV4LN8
DDzLHuxikboFpRmiYsH7SZqlaUQ/YPLA+TqhRAt0eE8dVZdEihuw+3Rqm2meZagc
biSkvIVJheH4hNS2hsop9792vVBYR0/VdpYrSoOMzN9QsaDeahuZoQzuqCZ9gKM9
Jt/OqJZArq4LXjF4DfRUBIqzDPA6FscpinzmY8SJIZgxmx5ZHFtK5eeRsUsHm0wD
YVSMgp/9xplS0Vrp4YGMR/eP6LRmDSTxaoHD3ixrhhUBJUD4x0popltjM8vNk+2Z
RY7BYaKPN39Qwr4xauAvSs98J3qBC2lKgyXJNin4qpH2TUjvO8HzZC1+nQUvNt2u
QqK/9h2ZjFMsW7h3SayIYy2f9/avxHqSWnmlM5aZM7TchfKS3eFBgqc3z8wgWcL2
ozr83wPot3Z8HweIwrFArj1XGdHGWsTQcSWiRHDWZeesm+71lq+11b+xYY+zbdrF
5SadhaGT2hqA0Wk0qM0QZoURZarQcPRqufymxOFU6+74mOkBYPH7HX61NlaHgF3M
aWaeZS+q2gfXzAXnjU6vxVwsyXjUe/mL1ml/VYkVneX+KJZ8LfczsOK+jMMAdgzH
FxNEufe2P6mwgtiziBoEq6NIHfxZKu7ZDN79L6XOtl2BALtHkTH4A3KZzvJFeWmZ
4Sm31GNzQWZht1igALEDgisCS173g9k285Qu1Bsy/0I+GKvRAVg628s+nJuu9fNx
Mz6+g4LG5fWgJ5WorhA3WxCl81ukhHPoTFGERlXvZ0HrZFsmGe1X+K1l2Y2FXEdO
6jVbV3b2Wjd3zM6CypchAlUz6E9eTg4vpJJhISbd0dZGdBYZPPHY+czGTLptkChU
3Gr+udx3VL4UjS+SrTulmTqDtNnj1Iz7F/4A5/lIvgjLTTDnre0FwspQMogE8UC0
nFqfrqGubSztKXIy5Arj6W447Ibj5IpR863NNNF7QbSCXddDA8vpjlT/PTSZGLLt
CgNLxJjMKQEYZi41R7XWNpUUF73I7faxJYxkpAUwRDmtrDnED1n8wzKw2ikJAeEH
nASPAajDf1YlVqARAk7TFAXGSRPVq4/Tn0oav8rnHT6ztp2cORY0nY6jap/qV2JP
5E4KG5hL5czsJeD6vIlXFBOeJBeXQeD+i5EwHdYvdxgOh9XFt/2pLhLRf9DsIo9P
EO8SCQrCjSj4GfoMbVmkG3l01CfD9mF2OJXgEKVgIF3ONw2gzpzWtDv/jAAoTZfU
0uCsAgvy3vOQZDoAsWQqcPa01uRyGT6sElQ3XrX68bX3UxXNpe+WG+LU9jFNaW1G
Gy3tCxTmsGnfvAuJ/sHh7zdO33/RlG0J2ehJ4RndEmMx7DTa+vM2YUG98VuXtkEv
vIWEzP0thmgPN6OH6AENimWVMzjhUO0dJGCC69cgPeFNIE30mTf/+VeZlwzb1Clk
OMLiYjhUnS0t3Emu+c7a/rorB+jyXMNFV4HgLDKtlzRIJJ5gr/BBAm0Pu7sFjJtV
zceW0VUk+/RJ/NVbTCsE05kyYo5LaDOmvPki0mZqS1GSnXTH+cPkY/tnUnvflP1P
qRVztr5JrD0yxKZLkb3sYL3jWz2cZDBMuloXNq6+TPabSZnRK8gI7QqiMMlGGlal
SnzrY6HEvous+IoABo3vy4Ss8qr7nTzPze2s3U8DfN/i4v81FWm3l2fwCRufvDRp
xqMSsJpAglGCu4zpQAmwBiNN4V1KQSh1bvBSIQ4ttASH6pnAXw5PdWj+fb4NMSOq
YYmBr4v/hcvCPhwSTE+ks4XsQ/XUThj1Y1D9Zi4XTatSZqbjHDwDkQEx4vREH+Br
aaIS0ce0soHAAmKudJt1myF17BdVN1+X2ev5sIvs7KeMjnq234ZV+3sxkvrhZ0st
wEtLaFhoTJOAcEZTxlSHEAHILObt0gDrY3mgdgGh0o8X9438aLwOtypf2x3L97KP
1PysDwcuxKaaMCKIxo4iwPh/+wOSj7ala9lcsnA6i9fAmtmgsQigAN2OK33vaIdB
cKRHRfsqzfwa32+LL59RX+HHbR5Zku9sHAxcvrx6QJDScDHjLSKrGDtMQtJjCgT0
zFhdsRAu83qp8o6f5xrTwan8OkwpAyF0GXUSGwzu6KqkkKGDX0WmIV+2I04KXUUg
0XJHv/EW+Y+yvKUb1JHaHcc/cQddmL9W3Lm6CH6F6ahfcMiLkUa/4UwdLIfFQ54w
EmB0/YFhWCLJuZGvpfW1wx6Uw8cOek0GzmMCBqHgOA0arllRO9rhJLctknKBlp0+
8FwwotNKMrXN8p2Cjr+SXQFMS+FcXuArCLn79sR1/RCB+QYUiDzujOI9cb0uMrF5
9WnrCJgqSQANYRG+5wOzCteYqOEG2zZoywnYze1aN0ZlOPNBeO2WeHGLpF4ker8I
Mp/6fMxrTP13mWzdicW0BA6VFpuYPaLsDTeH9VuiW4JB3CXhCYmDaodWZhKczVYy
QqpS2moM9hs+Rsd9Ubg+IrFhRNW+wtp/cK1OCeolnZbPHHhN8RDYI9YyTTpHzduW
TCLvltr3rbDWV+JS22usddnRsCVL3YjKRal6HqF0TFni1MhJR+AE9IaKBFQ+6cDg
aiGMn02JuHaqaLZabG9Nv9YkRFycrKzjNVXkzrK7hdkEHQefVxU3FF+pDaihx+IK
cqlSpvPxDDoTwM7XIUVpsy7H3CFV0cuQRrfZCopZ/Zh70GYxtcnam4T/CVmMTPff
u/RNki8WvrqOfiisNWFc8E+wgYUxByPGftkVhfbdob2RR4t6cuUk+aves15neTf3
DCvJ7rZiiMR9jqos7gVb64zGB7NkSPprgj0/RupCeZnBMyvY50NkRCa5zASLi7Ac
/9DhjbF+4d9xmBLn2IkuPBi0B+m6cDxXC24j0nyBPiD6fneFnkkahu2F8+S79P+n
kedNmTy6kueYUiYYu/zJOav/kjlL2H/J+Hvxoau+Zyh8ODPVdTZfO1n/NOTytOgV
9LlgpZ9C188R1ySP8xunDd1+mZ6ynUhkbeFXGPyDCINu9JVXAIIaxxTT6XAwlYVL
ZPLMtBsoR5r8QYnsyR4h5NB4StHX50P8QSf8UexuY/yJ4vPSD60hNGlV3EMLengc
JCHM4vlUKf7gSQ9RR0KuHMDh+HCgxBIUpxPq5tLk/mRDMC/JP7KL1czmFwbwzjwe
VEFmAHtkpt5uWhZMKSfibA2lscSellrloW/y7JCS3xnVsVpj6c1pHJejMd0mfY+W
4WfgtTsyom23VBHitmHH8HUOtg81XxseReIuIGeuFz/unG+QIJup763PgikOpbE9
2b/KR5gqL2+xW4gZuesPCdSdXDV5X1Wire+JF7qg7Ew3WUxneOAFe2S3xfVBnWI1
6q+DfRbd9AK4y3AtFbtmRhylcjQ3rurDxU513l2SlpygpbWbezrzfuetYqxuji5F
298YTfIoz2pxw9x+utkkU0xyxfZcKUIPpYCpFLsLZKNbVfd2YW+SshrWG7UdRLXH
OjsCnpmnw7bxFg3l2VyMCaM7oxLKAm7LKxeXInJfmvpR5YrZ7I3nt7SCR+hDLFu4
yJzD5lZsDbgrZpJRXMrftiiEApUOtlzXX/1njIJEIOrXUiWqYsIbG5m7tJobJL3Z
CKzMull2pzqIfbWn67vNhm0v2VbyF9dnsepboFFd7CmYQmYSXqt+XNyj+R1bG09s
DuGC8S7D/FfUw9SUw0q/ACv4ZIYpQbpHBnPGaaeF75NeHOSXOEWJ1rH+u0XFY+a0
wnMCNzfJCPCEhUIXWtmdWVz0t1Ffy9vSBhiqpyuksW9Mc2wuj5UWgNolBzBHdiok
c01B4DCVqJe8XfXNUh+ejUYier3XeEb3qn/RwM/qMkwdnC4RolPLdrWDWPmUhHc9
bavwSSwvSWRiDCEiSAuC4pPWu1zT5x17SZ0b5nGBV4DThgVyeuH+ELsCYnPMSlnU
btq4uVGyKrn0Eav9ApqYJZqzY8CsSit1qmsPYBBSbYXNlC9ERaXElRLfIbLngmNf
0+Q7n4Tp81LrSkmqGgI5KFZ0JK+MKqL8lXeetrUt1uxC0JU145OKjlwr/oROUYBH
5aHDZZOwk48pYHzDB1ggME/izN/a3Zo34nckNI0W9oke2wgN2niC7/nj/Z1qdQx/
OsNO0yK/OelTL5PdgL+E0cp//Uwb+lnV2CRqPkFcbNu0RFXfPghRgZrvSC+/f1/H
WgEzJIQbBeCKARqS5d8e9IZVCUsDUkkaIn6fTDVXRPZHh+fcYAUrVbiogU/u8PrV
oTqRn554hwDU3ByuUuNvI9vuCr1xToL1hfzuJVeFKwt4sH1Lu0evoqt7Pxpw4yXL
/wa6Lm3EPbJMYAsFQcxvbAY8+j9+2CjVbtEYlpnPzPwkiCeWdrf0hQfe7oltY6ki
LNQxOMVYhsKHo9dfgc3RdEmh2MKPyIrxPRyjv+iXDbjW5+fgutYzqu7Zwk2tN/y+
sxnKWAQmruRbgVAvKYPTBOF61K6sciXc4a2RjH53q0/p49Jz8JqBFfVTdhHxRJ5r
+1QfaQMh+Ag/92OOgl5Xh8hv2sCWE8ACwuol1Hq9Ao0qnuy31QypsJT4v6JzQHjB
oOY3cNNCk8Upf0D7w74bH71DJImQBTeeYu/wXDja2WBj5REHCTk/PfbgsZSsB3X7
vxvF1/AYejMZtQQll3Roe5gc1I043YWo0CNEX73hr4IumKLgBk2LEzm4IJ/pxhBy
8ryUM53fglK3TJeos++7UJxW3zKw1raLZfCYzqdXTlhYybjPRcVZY5Po+MHIGR0Z
mi1EloNvf6/wVMb2SNo+o/08waCIDQ9v+ATI1qU4H3fUAFuzei2ChB3XstLrqGoa
DPEzxpWfR7viMb5j6ceaFMKCt4h45voB9rBNpBDlFcLPlg1IlVxBQ7ZLp1KkclGT
YwVNLI9a8x8B2z6y7/hZMoK7OmkgiAe1+I7YD/VTdvW9aADsv6ZjnPlguPj+55vN
jG1bouCdIeSi7vA9dwf1m8f/3wR8aI8vihOSo2HlRR1JAPRS9LrQ2q/hwEizrAnv
ifskDAHWtLdmCWbDXfxpwZoS/ktDnTGmd0p8pk0l1TRa2cGgb/hwuc1iLZ1g+4DT
ybmsLICQeFbTmCE3CEiCTBo8tUQvXqWS7YZjZo0+N4TbTx/sCfpiCksRFb2CD4kO
IVWi2vIc4WBlkmAxQLEwlms9qx/DwNqdGZIpdeBRqoiJPB/VKshf5pN5BG0lMUz8
RtHCDlhHuTIiKrOlgDgbAP/Zhu1Id94wa+ZzQHVtiONP41prZWsgXb8UCeZeP3Vq
43SsQaPlgS3Sf1e1FXyWGJeEgDu/VYtnM7Vl2MZ7WIeCsFD4xWheSCVUEEq0XMMA
38kRqCnHvvkl6maRfCHDHWczPrwdFxaez5OU6kxYG2lAnY7sMrs43xYDgRcPavE5
fTw/qnn8XFFyWQW/z+HjzewJf4zlIckGu4biJVsd3IzaT8feIOCnLtXU6aqihMPg
6L7zR7lMkQNEc6v9MhfjwaaaoHLXSxVICNMWhMY3MtLITPyamfUMnO7q5KUN/UvW
1Z4IGsDWVtFdhaSRb36AtwX+x9c/k+86OfwdLDglMcIu73tiEaqzDG0EOFqKXf9a
HEAb7WaV+FNOAO5BSy9yinrwRRXeoT/zvmpLtxG7fETAJOCjc40pLMY4iQdy9A53
Se5C1usK9VeqijZzagE+iWbAhuwvr6XrsBcU31a7mfpihEde7qowDimTV49fRFYn
mczrkxAnerNEooJNy3q9zKUpfbCPxQg9WVv6wMXTzACeHXyiYb/5B9IN2GS9tzeH
wGWGt4T+6i3eTf4s+j1gSAhagIGYre9BsF0UgmrP6WyMB2KuZZayv2w9cFDDP7u0
Tn3DjB6GA3pozhPILsQm64ulvLgjk48f+5C3VZ5OU9eGbDBP/EZ/OpNrptZr5Zdz
Xrt+CXa8SimyHoQjPlMSfqvjBIpl0cJb61hxWjZtSDU9lNe39G8ze614BCkpJmVW
/VMSEIYFBXDrglWyyuvTQ6bfiVbAHtoWrXN0d6EUKCWbfD9VxJCtSnzbHHM9MdOv
SRA9HmrqA2EnyTr/95rCoPFPLfbeTGWtOU+suBbIFJBd7c7JslluUMiFo+KWJurg
Ds0xccn82dxUwVpAD6HA3Jqmp8A9UnVvoNk3HT3juVR9uLXYbi8ooAlSjYLuOYDB
ZhJ1vQtb0HRzTkXmnUGtQ0ELrr/hu2nYagyNZMynuglblWXf8sDvZJnp7B6pZtvq
xQVNGs0E1iLoM/ubkMbbpvLFg2iyxUd6DyADR5kNGLtnFhCU3tJsawcjvjSTUekc
wFeRCEGfdryNKrz1+rI8S3To402lLyJ8rj3GJ9+B9BgBUzzYndP695zwn353OU8B
gDbGeRhFPMl5YcYbgY9blTuJAlESKCL97DWWBBjBVoHeDg+Ua5C+jtQVkF5VXDpq
kKVShZdQwZwXpNSBfkRuFARO+nuRiivfwvnBX8u4BTrZTvb76ZFFtlZFYipEwZ9q
wQgivHdumeaDgIk7zb/bXtq9mdLdL/kLAdFvfr0jPOWi59lHfxTxVKCe3yquJhC7
HCuf+AKoJbtZ6j9RmrUTTYRnGq8HFqnBQM76vFoDUVQowDS+vqE5m0oeBfmiU14t
x86iPp/dcztiqo4QpZJw1NIN6x/HFbHzdg82co66hap75+4pg6HybW2nQIeQ3UVu
o0PKjFsU++0Ez18+96he0n2o9yc1PXC29yGPpcVG9jRcrr3UE9aZuT+g7by1wIth
Em7OjUVVGN3Z+yTiUhxvvFTssJwAJK7je7LwwcW4/qOMK82+ma3hbQFyjbkvp8z1
sg1SoebE+ggNvtuXGIF4VpaEWFi7Tv0cYpTvohb0GVLifb3e5/icMV3o57svODHA
fEij4vDJVc+9X2qAFeYWpdwgbr7offPHnubYiVoqDuCqIIcHzapBxzGC29IRm/4Q
Z55WR9TYNCbeY1j4ZagTyXpDfVdKRQWjctHKTyqOBo9rWHhbAMeetuDUgal57nPA
dYrZTS3hT3Vy8nQ0Bo/VygHxefgJlIUvHhb4gptUQ3QRjKZ1jCKLL0G0x2kgy/kI
Pybj31R0wDS0IGRb6W2O92J5ZZkHtBrFmOKB2P0hY9ksO7UZjaLSZYozh0OxlJf9
5CKG0n960a2qQWZUYrtSNjuCjCFKVInWf/LjwdkYKi89fYSyaPl2P5BKZCVFqEP8
RFzujZLYDUjTpgXQhE39mOYTCUdpUprPmrBH8rJgjA9VbrFk9drYfQ9l49oRNTsx
kjPQurp4+9tQdBWtUC7kQ1NdgMlfO9G3ZeclqDa3kZt7V3qGYKLZ20aHOrZhaeXr
GpcnFguW8Mww7Ef4uIb6qoNH9UOpr5gWRcUgn5jQMjG633i7/mI5b6Rx6c9DOvPB
A8JsIZUO0RFevhnk0SO6SS3Gc//gl4wrIYcOiyBLILkxAt1+U2pAjOnCo6tGv8ff
qyPM64ASloxwMkeUgBajZvw7Bji6KHrGS46u5R6Et4GSoPNSrKtlbI4npOrkqTc4
QEu8K+E3xam4m9KU5PxVYHtPP3vye6hpDu9c43ZvA6EeyPwPXTtjdSBaWlVsyaSO
jSZn8E6oMn4vMhefnlWEXuvWYcxmpjqzjUSvbgTQKAqaZO+jxOitGRT40dpQTqD2
6lN9XYW1FZxvANuY+8/iBNXKkhVR4mdoGvK/wBP+rTy0e/tOCLZk3JcVnbrKdtaY
kIUxkYG0kiOWUIdoxj7qy5h1cdIJ1vuUgae2OankLNaGEiIjGJxSbcRfOIMollcU
N8su+GORONUnA2wrWaXqu2X4wiVFwKL3qHv4B0ZXRaynD2wtGdKWQ905WYa4kqO3
BGc/UKzeEyr3nURZQm0KTrLuTHBmKyncXGVuN5C6p+Yt4qg6Ro3dFEZWnVRCfdW5
HdX2XtwVbnIiO1k538VEeZ9mBIE1AJvLpH3cBagR2+3gV8MVGw9CJ3XcR5rARcHB
KogCaTH4Z3zthQps6xnxmZNx9Vf3bNRvR/cALEXhCr6yXVuSo6gNEPOLPFXLVgtD
xTZSDMeT0nTMCoD7xLxA1KOJB7YvU2rfNPtk52pnuddZwo2R6jUpv5XGxK0/7Awa
nEJn0Jww2ZIMT/ul4Uwa2d3gfAgmX+HZyCjNLoGdYH/9tKXWDoX0iE90iFddsMhh
3s50J9XotwscP4kdWYANNe1RFo4XOqfA5AN2BlD9WnwNtQOMmJybG/WRt4O6EMSB
VTnjkERs+zOWouZhiIgaAkrKTH8L2x9qy6PYjo2Bf98rjNZXasg7Ez4nnkAMsBAj
ViJLrAJRvyxLPP8kPb6EcRLfuVY4KeNPRqHU5Cc6oc+teFKdr6Y0WEQ4cTLP8m8e
axfL7ICdFV/ljyISRffgnSeEzL34Ha4p024Ejz4i0kAZgbD2bMMP49iZ+GMqCiqA
sheTC3MFXOe3ci9EsxBiJ68ya7hFnt5d5Jzdcj8OF6TjYVl4uue/7c85Xd/TvYjy
Wb7WkeVfnU8HeYHinqTH+w1UlrIGLIAcxqJrfmswk4U1O8JTd+Qe3Cdtxs8Yr8t+
BAEuh6N2QDgasq6cxwni+xZ1v1o/mnjIZiybsYz70N/3DZAyfB/nFs0I1v1bnZAz
PYsueoe7M1g5Py+odcqhkdSMlSqnfHy4W5N0sw75qgZoQ8YJJawtgrFwNrJeaVn8
HiiZksAmwgXjA3oboktNlaPsK86vgDBal71ySlzLVAPSFQ/s4zzUIzwFzyFDKel6
JpOldh8FNYHbuTgCjgI0/1NvBNlR2uKDJJ25+y9+EDV+5z0bbnejH7kluX6psyKz
pDEuQnpKNZH+B+q0seWXRS/O2CASokc7Xr2xAZKnpw6rMAfS7pqc1Ygxa9da/czn
lqQQrPqmTZ9niIThp07688Pp5KUHbAeocBm6kGmpL+Pj9tuFQp9T4mFcEtSszoAP
4GVy9DVkjyFPgcvmKhjoSo9Z8D8tDzyrVIB+/2iwydc4/mUnA8cOC2tEA3bH7zQM
9KLzwwd0H+tc1sFOz3KFo34UKrJtZm/qKYBhB1SUSO90GxQcPilwCSOg/OViCfcr
yMT4w62tWzqZ8qW0nRzggGqhpjWjXoK1TeBgWCAU3zW3Hr8iY2Zr8WxkmsxM42ps
sL/oPt3aWBLYZD/4FIcu8WbErjwuFqP70NIQKEsv9xICNuw/ehMvPaiTDzof3312
BQyCF+RfoYDweIdGLIWDY3CCJkj/vNXTiX7/XtRx4cI8CFTbKnwgoCyQFpmGPl1P
ebCFze0VKiEu1AMqpJr4xx8OShmRcFnMeyaR+TSRyIqwXiJEvENtq9Ls+gwke0HI
Fjx7LufzuCr++3fgNLClYtiHRBWN5cb2Hc9jJ1qZYT3rtpak5weUSGdqZSnp78ph
IOOK1d7GS2re5p90iN8S8uJa5YivGUVvhI4DJAiSBWRjj+GwnlgnNfHObo8gc81x
x0abbn4IW4gilSespHz5E45ENrb6Pfl7o6IHlNyjUJE1qZ2oX/vMgxok5K50pafH
gSi+erWa5mm9ZPD0QzAtLO2HQE3W34mvxCpHrMThScB+/lnB0TRkARfI3TpCwkgA
yexxb0jFuTBLYJFCnf2O453xPwoVJlsurImgjHPLDo0s3qgtTRldCZEzrSNklMD0
5d5vemC12KF9x24IGGwPox6ZbZJaiePRDbLG8zho2hk++dqE6rAmPF2Tn66E1fKh
Nw1SvzAK8njUt/a6sqA1/6NLfs5yCvlM4ODUU1YHivR0NuQ0TlejMtl8J/uD6nDt
TCBxlAhPSFcdsDk/UzqQPIpbx7wlkv0Ty9NwvC3sHkMrQ2AdU2JX7r0kU7s6bRXM
NfHFl/QPrR5LmKiEg6eVGsM1YJooTFXdipijNkhHxxqVBBdelEjs66q5IRO7zvhG
1xrVI88f4Qo8XiKt/aC3408uCzdVoC8PWGoTeIiJQ621Df58SsmXpg69grgYsiIY
u9a0O5/KxJo5qajBWdNQ2z0JQ6bIwuQpqky3qdxp8ehubUZE7LJz5WbOGFeo9pEp
1AetK21/LoqXqIaYWiVkgVdP1FIIfAtxHxpJ7dyekNs4UDeDhMc+htrP9eMZQB36
4l7hBVFjmaiCyRtiODkCa/Uvm3R4DwzvQaYkPTqV7TEk7ocyCxeuDD0yy5sU+QSn
PIKCgGct4lW1DakY5p+Z3qXIEsA+n9BJ7ZRH67eFzBITKRr8yVEF8163fzrdSvrT
Ln3YLso6BTYMQMlKB5rYJAIqBqDIf3WRoW6gSZUGlG+9Onjf3YK4Gw/37ZKc72Pn
/DZdz7E+e/uWRU4aL2+v5MyK7k7n8OiW0YU3mXBrxaM4R8O6eoMsQrqgdObYjj9k
kSLqsboFDL+6TVbs77hSVFnMPJc0Cb2MTA+18d2XaQFpw1nmpFoUK4gnnorZxzcn
yLBlxjByWV250olYg6vHO3++3daCg87KXcy/zLEjHfnD2QIiF/XXTFUQZ6gT+/oG
AW7CdK9Il60TmlZwPGQOm80u4bFFKSI63GQ124l2uv7haLr5Dm9yRgS/YmHpc9QK
oZ01oEsv9vKmeNPNLqelP2oz3SBEqTtJ8iKevHK0JOJcM3wBvGrZsWUqGQS2OAQo
/3Q/0CqgcZjovhqhMyJrpeVnxi1sBUO6KjI/j3NM8kWeaQfu2EPTu9a2MelluvfA
aLPzw0VE7P1V3MxMOwxRGe5JJ3WfskJjMP8tStUbvetTu4VbdqnqrIRnyysQ0Qmq
u0V0j1Cc+qnVRZZRM7EVVjy9w7V4liCJ+AlDrL7MOFz1oTerY43GjX6JOEFATHoy
cSI6Ja0c4pCorfVKGWxAdjpc1EVd3CtZW5+sVRFs+bU8jXf7NNXKoXsYu6wgDiyj
CaQPqe8HF17XBJxkXG5zd7gcN5XleushmQlVW/Iu9LkkHOCl2+PhyfJuBHy1Lza4
i2BaP9IAbx5xkFaroenxcx9ufUsoK4K4iMOLE4UwqQx2VFexLWSvryzzdomVWaP1
DIMH1YQn+dx9QtR6zqmaogbghmY8amXFPLpP6AMFM71wUjdgNYLgFJ9Om2LMpxFJ
76ywNTQDV8Hlg/Yfvuy4Jcla26yzwauW7QHSzQSCTJAhTWQoiqdfYoRX1yBQlZ3N
7L9/eSBOWRLE1OM9TtCRu96sIHaAA3XTWINs09pLDB2HO6FpXg7nUcS8Un2n2La6
TfJYI2XaWDtWNIfzOxs6C+kaLC0JFCuvJp9i/CrV6X9Lgvt7QQepev3M1VcUhv0b
8kqWycyjKgle3Rf0rfDEJNjajTMY2AJdCHdEf4FpvEOx8Hk57Nqt2NvNFFxNC3Aq
mCU581Lsq3fN9TO2hKeZ028RMkm0vB90h3xcJnAgoVBnbsNNQmp4H/fIuw3C5vpm
e2qMJJMZF8QjyLbuR3HhCa2ql6DeyUmX+xf4qIcCCpLHtykx+9M8lD1paXeWaQXc
3/iuoDD02hdMsZXP4+XH8merHWup7m5NX5B7dAJP3TaPPbVChS3uWJ2ZCFWiDFMc
Z0GtI5g5/r3D1FMXuGGvEGVxm07CJqjJz3EmCRWTuV/tv7aNJa+mHpg3VJgq72Ek
N6GQPX91jaj65jBx/LKwceZ5yX7xn9Pe0+NNV9d56wwl9/IZFgrTciW5BtbzUEkn
kuThib+H2gZ6VMvKVJvaGB9+ZNr+d1t2mm592N2GaQSsqS55G9zGkT6iP0qsEjN4
51Ce1vM6rt4FqAc3X5wSM3Os/xcvrQex+6FHALQud+hw3Pk8TZs/yXRDKKvLWire
GGQqq8Z4oQ94nNdm3WWLp+gTeLCuMjEgpEekP2/Pz5JslwixRb2FIEKnw1UGHH3B
IlChW5erQA5YkyPOLmI7YpoifA2EdlBPgl5P3PlTYBCHu53hXEdNk1/7narINt/V
UlBTgh51qvm88LleuSo9yK+7S6nHO2Pkn7HEyOiwaGQfjSwd5IEPCFgv9exg6VLU
PwaMm17TxlJ8MsrAPuQGqeqX4KWxhVJiC+EY7e17uFoWDZBIP9ct/XxPNZVxqG+Y
mJPtdv3DgjrOZSTPhMbr6scrK2ZQAbgF1YxjT+HjQRFacxW5FyOq7SBbTb4N5CDy
kbIwUMPRzWtvmaYIkWek7aURufD0M3kv3P7Ui/00xtrb/1lVzTvHO8wM1cmFO3TF
Jfk4xwQDN3n23ZRVH+iE/K7RQBvLkltyfeCNDECwO++TuZLV2v3/7IRcgJC8MxmK
X6TOw4mL1zD3PCFp1q6eNpBIJSVAllV3eU5dZ4XnJjOAcHUDK5xAPNW+bi1QZS6+
VqK9Q7fjxrvOTtcvnzhE3VQXP0ZwVmTXbhcrSNDMLdhhSU97ZP9+/IxfuUbXnPLr
NPXzC0XjhfLhs+zSTPSyPlXGbwYFa6Bp7TZW7KrNn5DcveT12cz7iZDXp6v5NkRm
UevEnK0XMBqwjyjnBfA42RjjFvezCn/m9GP+U5eyJEmHbMaeeQUlSijPmWU4PM3x
Fc4FGsW0aOfFefhpomzmW0FWuC4fbuRgK9zwHnTpnCHapY4kHcuSZWVqSIHPMD1c
WhlZk+fjTulZQc+qZDNi2MKt8MqL9Jskv7Hesyt1emiOotSlqvT2PPjsm7s/L/cV
4YzuDFz9r96cGMb5ee0XZa16NEa6kx8LazvK6Km/tR1MA3dxzoeu0nQUUJpkE8ms
FOVTV6FyrvQlIbq59dYMKpxA+atsAeA9bCjrbmmzlWshK6DvY5+Eezv49k/m+7an
MV1u8zrY5Jrdy/oArkiV9XQ9QChNjP1OD88gfLOg/cqikuYv5QszAu6EpmaaJ2aM
jRZFxi6kiz8RGetGK9RECjDdc/qnjksdzZ+o1YjTzga7DLObZrAjqem9l5WeZ1Q0
kbPrPFxh9Lxrm9mh4LqCbjv4jzQ2pLvu136QBVMeU5HckuUlCORXOL7Y0w4hKlI0
ND97dGF7fAHVqlMZmyPdmuNJkBBaCoFw2uFjVQGA383mEdy4S2gj0wxO/I3m7uyh
L/Z6dmlSBBVQevItUuGFXR4QX6M0obC86MvjzcJYIqaS/vB4bfRGkRl4rWQItPkc
EZdUuX0SUA1TOUU7YxPWF0v23Otz7kEIhwPMh73/vS9NjK5EgZFBYrzH9DIO7wqP
DEtBOz4KCRbJl8RHU7JmM8gIWtiP6SeLi2I7m9qrmFKzV7v94tm2ObMltplPHYoK
J3h29mWdxRRowXYH0zSZxhUWgrMYJDuoTV3ID58A1nqfoiBqXWda7TZ+4N9viN0z
K7LjSbR5GvWfTxVCT5gpFeiMV1D29NLs91ih+Q/KkMGbaeOwG+lOY3mqOwpNWiYr
siz0zQpkQyqBoWhgyplTKelKMBErsmVw/QRfoOx1jubULz+iQha9SGIMUCS8nbLW
CSWKERuKYbJ4RF2Wt+qffzBrM+1AVPnSVUhrZZHIPmPvzkPWpYwcLE0T8mpIiDnO
7pLYJJUfD8pF3lxkfjrX98SwRbRUUHNoJC9gItZZ33nEmjMn4xZxjp7D4afnKbEN
/6Zq9L1v72Eq8J4bynVplSSBFlB77rEqi5x8HokqDpcBmsOky+9RGDzjCCc8YxsG
S88HOwJKQctnRRhh+u+E/eniX0MFRN99BPzmcVYzBQ0FSBlm+X1XZUbaZsQ+zpNt
uvxncyBEIvNaoniO8ByJSYgzlqXAwkeEbyNF9TPUe7aW0Iz5un1CtlUVYS135rXy
F8rzTIhDLBVusXFYKv4GoU4eoG2FUSpTIY6fETD1ZL3lfz3U//+hWE3JP3w0ukUr
fle2Zl81TyINOo16WyNcg0kDtxUQv1vlsiWcXtB7b/y1BWkwj4fkd4azZncT8Nxl
lRvrkYzENsg+IfvdWTABUR6D2+EBEND8OQVz67aeAofYSGzMpxyceDVd9gAeEENc
UYTc2wBe+YmSvGWRGQ1aKWPJrHJASayATZfCOtbb/dw6y09aSU685+LYjr1dn1Ww
ejydPypmIkbhT5F3wcYdkMibQYEzAZ2mQlAxY/SOfGhMeTIh8zHwSZ9T5tK64Zkt
RAjcAqWaJAtywSCYEmZIhqoJsHUoVB4OwFuHLb2YzFUGiljdlOX+LGUl3FZE1/oe
yf9yO0WLK5R7d5/ZAe7tc4/H2a2gdG0o7uQKaX2V8v0XzYYRg8/k4+dEkfvoS8hc
pxNEtjqSbSAgnHsFVuMRBv8ZcXoOPsH4ZSbCxgL1NMFWNo/b+zeH7zDQtBBmBEje
5fpM1JyFWgn8mKyiuOnogBwlb7/r6ZKl/YNwUkbTY4pJ3+EBbg8AZ0OP3gFDFLTV
fxC0fJa70o3FqQrih8U/s7HhBeP8eKMKI3FxrztmHYXEcEu3RYEgykQu8zdzF0xU
R9vfhRsUj1MtI2wGzKVzPFTobVwGEi7F72nfSWn+TYGlaYrvHJZa89Oe/ivZnAen
PwR0aM+pdqFgFCyzh23TvSTSn5YvMaUFOZ1aeNA197wVeCoG06nP2AuDITHEzbxK
4bKcYqY7+j3S1SIRF9R0mbPRM9Xn85RuUaYaE910+P+3MnfKGULmPzriGTCVqjxi
WyxOTjkOiI3XAA3ssCiyU4/ysWwaMHwlpmgrPql3j9XOB0XkcqwfsnfoSwZP5E5r
xgeoEFLD6wbhL3TmuP4eVJnBbcxWg/fEoIByswpYtDuyTBBsCgE1hcRmssivGKYq
wVI5Fp9vMfMFl41R9D9wCOW6gCTHVqOSpp6cCO4D99sxbfyBwU4SLQ7JwXNjQ5oi
hsscpvDcgJ/gOQo1AjQU4l307eECb6FIC82txQtvmAevCBRCYWO7QcmSo1bh4+pN
UjNUMlW/CUDVrEeWQrr4elwLyopC9YGyZZe3hxyepZjebK+P9iDl8mqNAmwTMpYF
t3yAEj0hFixiWGPM5n4aGDxDw/CYdJrC9fsQ0++rlHm0Oq2NL+lHA15XJgnnTWUs
UMi5csAytNCLkGjdgKNJNjuTPYIencUFDK/hI90uKJ6ePmlyDy6KnZ2G3yX6uhQh
DuN7qecs/anbrLa45SMJ7Fc/UXv/qedPSnT+NZnVM8eIrGMknsK1hGvl59vX5MFa
gYCGgNQFaxGXSeIzsL2ifGAieJw0gDX3LbuMQFBuBMoHay71Cd6lLVIczPz5PiRG
ry3tZY1abCYwVFWOGGTp+hwUxGnNJ3oOJXOQgTtYWupB4QoIovxEkuohYhKa/pKg
q/ARBPSBNrA4aZvWSs/ASU+RsiM7ooj7kRTb6tyMqmHeHrSYnDXOdnIygZpNZ2WP
7z7jDek+NfRFZA3tfoFK2ECJRrsI2vluwkQhiYRkLwyGl36P6uQqkfnXDiREiOK4
S0X7ya8QoUDdIbTshv2F/T/lrads95KKjDvxzvZ0hNK9O7C5O3jn/OORQQxXf1Zn
N/Z0FB/B0uEoV2cM0CMeTSrBPdsBefppzrO+Ujgo5ukEm7LArH/omLfYphx7DxSk
ROu7GeR9YYneVf+HXjujPMXn3Ai5VH5jFQfrraTPB0uuUdToHIw5BUSLUxrA24su
MwAI0q2EXef0C32r/9CFktrNy+12VX8DAAgOQ8ysJ+2QTIbhSasnkCNSdgTOIJCd
mA9xpCuQb8L5AnDguLMxb3EiHCDCK51HOp4pE5UfaZ7NXO0l2WVenWnTslgncwK1
pJF3bTzvMOakG0n4BTdfqQoT83Kki968MCnxSIHp4NlW/0dbYBWcdxrFi1N6oYzX
6x/U+2LqzpgIsivr/I1XTE02bAARwK/1dXZnIkXLv38SjB9p0aPSaIgsffiIy+9Y
Qa6TE5y9JTykq0kvj1hWCu/j4i9rnAR3aKcds0bFNWZIXOFHj2DhkHlfFbjYONPH
aJBPIyeSgeKJ3NyNaKzSqc3/FKqPNCEAmCzTpty+hfQehalGIaxrpLB4fX8uAlEw
y9rqWti1C2xApAD0poxh6GtHqdEaLr/JvFBCNHnx1ifXcmjawgLSug/l+UbLocII
BRrVFCED/Eg3Dc3qS8Hg704/E+7kPNzITX70YVlPfAUqueUYd8tnrn9S4KS0MT0I
fgjNtr/Tgvavj5/VHMooHY9Prrm5j6vs4kgVj4lPsq1ANRr9uOkHxah6YNFTzuEu
RdZXeMp9j4bM1XvyFn0mbW4OK/Bu8kCcbsPh7754uDfCVL90G3m0O0jiYDYVshkZ
23axRYJQCAlR6nkp0Q0H5hVFhwA5HRCWRIPs70W+7/uWpW8V9/1VtbvVDtvH5pn6
JnQzSktammeTGqc7BMwsfGWPZI2mrMtSL0XODJ22iqYqfV1VImJvCQlU/Tiat5Nu
qrWqg6zoJFXN+IBG4yMnWkOazhMs6dTwbM+A6J9Ey5G5R8DJkYXeh8qSRiTI9X8d
Dr1ZQZYLxX5xkdJopjuU/5Mw5IRrVvh3WAui4HJ/naNLmtXfFHFR7hM6G0Ot9nFd
OpBYdhtrK21jT9wvVVCjJ/fSmOiKZp/szkyCOnu9+KCbzljH3YYRwYGAmbjGBSsT
TdsUHpjFpE8setkfKLXd7nuaLwQcP/C0xi9wVIvlPMgyB25PHJbVTNy3a2Txjcc3
WWs72q1BeayurrVy8H5u1ovq54mqgQYkplU/yCuPZB0JO7Kimo2RBrFB1lNCDdky
BaByqYVS5xSCGUJ5YRxvGnkLWFstNg8PCuliOgFEx4WbJF7O8Bl/VDKrZuYzGAin
n6sYxx11F/7h+emmzCbJovonVI+e/Gwrnt3VvQQL9wPi5nAzUl6BMceXb/THvTdA
6ACi9IsOcJdbv0Os4Hb8XH4YADGYdmty9Bp+gSpPAIaGgxUsRjcCmEdhv6EqQqhy
NtT4RhOlUpHu530N2SAGbw9VKHWrwFIL3ZPvO/gJ0Rfoj5Dr9ufBuUfPhAJMIZV8
p5W3wJNnRGLs+mlIfr8Iot/1tuYBuVj9/oa4QKnDT0DrBKmjyFePZqu0RY/zuH4D
xtlgpRoQ1nC1M4PR0avbLt1+UoM3ebR5EYAE2o90RfgR3J5BjBHdviczZTjhC2/e
A+8BnoZXEZad9aLk8+u0sf9I2eNlNIDsZecQ7abP+OUR9I+XD2klVSvH+NroDaqP
0D2jtArjOmlJQ5JJ2qLc01sRAyOdapDx2b/WXUVGQPZRtJnSKWA1mYTCljHxKJJo
QwsXV/Ze4lAUkCCOL1Sain9h+pyrGTlMYv1B+ljyG9xSIuuiiZNBcczFEjzucI2T
Y1xKHz8s0JOXcpsDtSlDj3n0wCsuawQ7v6h4vxzONeFuHYRhdZ8zWxzMhUVIgVMU
alsxBc9152m2VEQxk5w88IYRxr3MSFOWLzdL8tkT1TahkJ0KUlszG3T1JqVJe6RM
VCK1AOGwa2cLD8SNf5/p2ywFmypEhvs9vRMbnuI6Oxs01PevqdW5AWrf7+KBtvgV
TtfwDbyYvyqtSj35SVzlSHB9nqkxlPwL7erWEH61Ql38/wlx7WVRn8NDnYtziBg3
MyLr2SmoteZUsrtz2zfuFKnwTwKwn9Peio6ShsfzhgZEroB1Lw+jh1nNwlCifWoZ
lJP8iKZGfVkV3SNVoCu63fMEYMEpD3EsSWIB1wSBMq/bokarOf4evk+G9XwTqxFA
LWRMAcwTAE8v+Pu/rkzPJyP0ZjwLHxJEYGIQFkPQXWhJhJygZcUApV75RwLeBeZp
x9LaJmvarmrZ10tVAPOQjMpntXlLbQYUo9PTI9NGCN0X37RXv3le7TBet5Wd0k00
xKIeprWimSWCh1SxFlPXIWwVy6c8RwYibGNn+/K6l7cTddxWhYrbkZE/+KiOrdet
Robj0Ap+0i2D0wQU4f6gZJcwQf3CfwbsUw1eYnPzqPFhOR+33uCI1oL5Xu5qYgob
GK4GlzONcHfGq98O1j08KJQ7YT1KJPJDaZT4UluUdhPpGXSMYjZ6AYAZWtfj/A6V
qSwAXtAOR8YtgPU0Q/suQfG9zpBQaamnWdu8hquAnITVAEP8jzkZ7XqHQuHNB5he
OmAuRqe+RZOyqokfwJpVt3R4Bv3a58DP8mQp6x0aGs5a4rVv1OgqZOlxSA5blU1S
fkVfsMxRPvPRByCw7NdtVk3jSpqRDJLuMmJSx6xCAqZWPHlS3jZSx97f008lK9Sw
jCdzvdIEYioxywhj1VwWXSjz/DXSJwq0WdHXbwXYE4VD8DuGW+h+WG/icgJZdv+9
tKctTrxnwQXdManfa3zEAoPmpjT15uIBfHkVvcxnQ9mEC5ToWG/JBF23uEPZnmU1
PKrjhKM7xqlXgzvsP5EsP1HCzlsOgCNiehpAoc2/Cokw7TPZlLsl//0dp9Gt3mt/
iMT+lFre8pY4bjmBeWwEO5QpU/xDtQtzCuqXkHAZIGWhVn+YqajYt++iHBeWIiEy
srTgLJI/8VpcemuOm0roAnoUe2RGoAEiRt8CujmzPYOpuG8m+mYIXTjH0DZxHy0B
yXUcmuN/opYc3nVoYRd8X8ESFIhrZuhyuv465dSsHxzhseA5nBf2HjH0t6b1lfKA
1qWGnta5fXeNIYXrBPXnm1gOzUygfe4hj0X7Ulmc0RwbODxab0sFlWiNrZ78EBy9
MTjDoQ2mW0xViJ4Tizz3mROcsUhVP2dqTFWIz0s6vf78OSLov1UusM1oljjC4/Jb
mpG6G3IxvN+omOk9Oum+v8h1imdH3dkcVfornQxzRBqGu8QT0vXppDAMH+mRoAxu
hU6kseFEsp+V+i54T/iGTdI359VSI283Xi9qMWuF0T12t3C6fHsSpkUgyelOBbTh
ReEqTOGcI/DV5dQy8Rodp/CAP7Vm/f3hArBdtjeIoPyDnwGgxN/3p0cqh8vsXCfW
q65ExUaYta5Zh8P6WtRPvcFjUqgQ3cZfZeg5migGoHstdlIlB5knF+/FOwXCN5MU
rM+WfpwBjqP5ccuAFqJgLEU/o14M/Gq6UW+4cYO/MFDpCxs5CUPExHf/Eqx0VN5y
XjGVR2YbTaC3RUIAev2FAS6NY/wJCI/uFUZybAzgiVSP6webIP4dBMc8IEVKtqXJ
XDwUPPYVZSD6Vz+4dWTd4uUATX1p1BI6kshWpUaj3pEUONDzpKhW+RtetH0VtEQM
oj8HDaBe3HZWlzzdV4ZdHEtDhSB2/29CoUyCwN3rENSTwWX6E0fy2w3u4juVbQGz
dnWtmX3/+FtvmS/tDqWQmcKHFx2HUUAAZO2EsracT3P3Kok0ybriLjsMpthY7U/V
tNRgr2R/8+mvZmTBabBmeNZnQbO3ReHUeaGiBx/Bw3t6CtJzGb73Zu3fNcr0kswV
VWzWy782jIKtFZWys2K3iTO5XTGj5OTv2PkH86sTGpjZ5HZ9xFS8J9fCwrCl+Y7Q
auQQzgQ5tEp7xHFkTDgkxEvF4rajFq0nORvZBAIyFhooCHP17D8oaf3CCQO8khI0
xZTrQTxjVNZj0LvgD/Cf2t9uxE+Un/n9M3YsSKR2AI2REO2bE7ZYjBEd7BmTkEef
e/FBCOuaf6wDHePaj88ZTyRNtWPRUoh5BRUE7glq9G2tz92/ky78a9fC5CsCSuKa
urDQzyOkeTIapAwTwNJ/+TQg6W7K2X0iWoR5LifAxSeN7TBU8ozKQRoW1I9AcwM6
wJcN1H9JuEqV/CiWA4MNWOkZf5lzxNe4+g6ByqAtKvxGdj065ZSI+FLjqiYFVbqK
XX/A38VpED9fB7tSfp67KPdj2mnFBxIRVJ1NwYU3vDQ6oGlCTZ2EzeV3bV6NvM4s
AUwKg0BtKmASzApt0kWIUJjNpWgUD7hWLK1hnGDy/SsTIqnowKyeBs8B7fAYxsWB
dVB81BXLCIWhWK2Zm9g3MHcblJwcplLZaPjGVaGpkxB79iSMPgY5pNFHZTs77Fc6
SdMs6CQpM5yiXrdcCjemlvyIf/3Ai1/V1ufzw3vYcv2ABE17Abcr2CiAfrF5H25T
3E3rft3kAjRLKKg7VrlUVTlI0oNVqNfsnqIgd/uorZjsv1y5ONg+GHeKBkn2u7Lr
Hk4+porkxM0ijvrnOo7zvAA/11S/7ruyuKOan8DYuk3bZmI5cJAaa+fcrFbizrbE
J9zhduSDRC+Xov/61/Fkd9KEBxSUVkkDLlsoEOexRAx1mVYlXlqLusarx3eq6oOb
a9ZOJIlX3mlD1VIL0hECrZGGm5wdnoLNpyL2e6gPtMQhA6480dKGHqRJMhNpCd60
r0DfKnzIgS+vNxL4k8y12SgJS8O9Fy79KkhVxzj9KAeYLyf0LX9ZZOdxAvIEQcTh
Ct6962gNQGkeNXlaXGhzk2pAu3c+HkHaDzZHvuszogje8izBEgdjnVBqqKVyxsHq
/QnoVlUDTQG2AtFIZ2zvuaMXb0tyGpdkdX55qARNzeV345dWkVEofUON1cjlLHDV
1WaBVqXsu1nvp/aqsLB9Vif+eaBMjFfT7dRG9CFBbEqxzSd4n8FwsRmIE+rT8v9c
YbpagXIQ4HzczTaz43VpEq5qzGYE5b/kenlDWApsvLjQ4s4LuEDnYXE/Gr7XlWQx
WPMJfCJSoOEhuk2TtNpDWDRIwPmC2Ft4arGceKDcU9+j5cmiftLEAAK7vPkDPq7U
yt86cOPfOtBAQhQwJpWQ7Enb6vPOyMonnbzRrNIcavn1pO2J/4GVzmXE5R9OiNoo
omv8EMElR7si/v9dG8rzNgNYQxjQs+2F1HVv+MsYBbfcFRNVtyp8eXoH5oEklfJE
xK7ndCx+Ynbb2Jszbm/Nk5VVciwxN0UjC8uPylSig4awpNyTr+vXa0c4I1gfUufR
mjg/uBiUZFck7uUArlrr1MpLsNoTa7kfG3bmDqGysTtOyD98A6/Zj6HX45a44yg0
TiSK1/jLSq7yGo17oZQeQJ/cV9I4+kEtHbka3yaHk/6fb2+C14kLAttcNRvXbSKE
VOAX00JIk1mFET1gnQXY2BPrPcVQQ4jpD9IE1Gy0BIo97FnTG+MGAnc9cPzO+rdp
uOj0Kpdz9G3U9IhWMCbjGnZRIw+CoS9a7DZyq5x9bGUAn94LLczZNP5k9Nc0Ih3o
CiBaZVAesTX829FViN93JU04DzkCgyg43ic3g36mNAJKSRxqlRezNH9EIchrRIWk
JX8Av57zfkQb9klkaMeUb2XsnjoLpBnynzAGOBBuoXXBEfN9Rbd6RekzNoLT1yVV
o7wu7MEMMYz4Ea+F8K7CN9dzVHHlsMKgI4e8ahIpD6h8fv8ANrb4V9HqIABFaVk3
XCm2+8Aar4+WftBv99CldYeuvURq2kCBQ4/za3zQEWdgVvJtuzjlSjxE39Afa25M
qbYMQmdB2lQhzGhRmXvjFzZ8KMWg09Bww6sKILipKcniXTHnXv8CTdg4DAEzxTB6
OubIYAaTXCEbvI+l6DPrTH6sar+tubz2vdBt6pMpZDWhoLlucct0CkVwFUZG1ntl
jNiTPew3n0gnjpVENHIiIQu49woeap3xL4y1waoGVJSKa2E9Li6hSSzjrpZ/MZXW
g1LVg9AJFYel3kvG+4RAwcRkV2YD5bMvReuy3fakFKf1XarJg883TyModvz2+6rD
aQnpKJFlX5AP4TRLLMSLr1N8KdpVsSprjmYoUL7CFdPaYlYJkVk0JoOW0Le14RdA
8qWhs65I+64nuQod/aTAd5F9uQ02Syq/j0uL/WVMBE/pnd/m1hmZZ0SBtFP14vsY
Y7u4AZpyUlrU6XQcM514fPNmmfgfzqPrIC4GIK6nxW3ySZMVZ0iQuCIx24B4skAG
liAFrO/owXEaCYWiEHqZVHOlJE27629+9jqGWiLQ0v5NyNia9mP87tnHsnm8O+Ac
lcrEt8OBcoXwlpE9DomNcHTNqlL/51sTwKpCeCx3PzCwIvIEqG1+irAVT+qqfJCJ
X/BA7OhYxHyNE8xhY1QvPryEu2ScqMGnz9b2thrkq9vNZ0/K1ZjCSLmSxukxb7DY
eAS0wj+3Psn2V2jcVjeaVJXMCaTw4GFfJ4kGhZ0Kd7FGklut6X/XWj4BmbFV1fWF
7MQmLMURlTZo1ftEi9TYIGVorwOzHzFn9ofgUGLUj8DLNaaN2p3UhHQAwuShltLL
V5Ukz3Hvj8iGy1guS295bjatRmkHYJxgPCVgrddneH0VEmUD49qhMokShvr0raEQ
nMsjIwKMhJNkkASoAqJvfzOD513KRR2nChcgNZbzXB4MGH0rRlyXUeQRdtWMLWqR
CIdwXUoV0IdOiwx1C6EyLT+/rX0vBBDz+/VTm+d+YQ5MGffK99bdgg2v2qAGW3vv
lKT/1dG7+56JpYlu+l3ymT14USq1HBwE0xFs/PesfYLYYqnGgRj3Dz+L+XxE7hu3
GY39OHb051PO66pmm1IBajw1Uf0EECBtCh3vOrKoSfjvc+gl3UVwlqQNo+Mu9M9o
dNoJw89jreLKO/oOCtBYp5iyOfw0tvzzubOSLZZWX1WQlW98aTKtVbaQjVB5OlCm
us0qqSx1moVAeRTzas6hMc/16K5pRc3g/I9kfQW/8jl7bDTeL5xJsunV8GTFtCan
rIFn1wfTppsAQaYEmlKt9uc9+7s+D71b+cAVuxFNxavmpS6ybry6TO9fTJt3h1Y/
RWfeBWzaXjfDYC8PGgEdXwYYmNvbVSUCYJ9uZ0evSeJTPI2SXQ5fHT2UmDsrD6X3
pZ8HyBnKLSIUgr39Foa+8Aqi0YOeeNk/uoSibR6ldUssmBHiLfuUbf+Jm/v+WJRZ
a3O4fveVz/4de45O6BPdSwuzKK0d1czteBixudji3fYNhfyZLwkA9Z52ZAaEmzBn
NzEiTFcS3OT39x7DeG/tqcBzd6oXpa+7u9l9PRbYsmhT80jLDKQYAxiAtGB354pI
Q9t57jtoW8vuHeEU8cnT9Px5/1TonXH2eDvqai7MVtTy6dlp0r+dS+xkjqSB9Cz1
2xrQ9w+IKIkXM4PWB2mO2c/Zr2EvZzlU6a+WKBojRtwOLIeJieqjUYkk1gTu4OyN
JAgAoOEFyXVdYaxKftRA5mGnpxUhlzpArM+wOfzR9NswHY0QVn8AcuM6IaSk1e6q
2JlzxvWZ/PBdCJHzGPLgx1lkoA92BawrgCr25/nQYzshxUvdbBHMzP6GfumUP60U
YtzfDh/1OtPVigvux1fGMPzVJrlQXJkIntmWJDmQFvqSxIyOrK5nUwn5HsR7TxkY
kuhVdohRxDCNNzo9qB7WxZr5QAd/hB30aXah3ASInQyKlavjFWGKhsSH7TP5L05f
JeoN49+ftPFtCfIHPK8+JfQCFmUEH1upEhPtgyBczUuEhoxuUoHKqGXLD+sfIfzn
Ui+hf7i7BI+YcHoe1nGzt/Ms7HhdNepu+3uiMpbHEeJGTBkq+BqkWmhh+0oIkM38
erUTfI0S9dEvDZRjk/qcdKWQ0GlJHROuzO8dbDXhBh4imRQ+OYk6c8C3bbWw5gI5
gL2HaQcPLF2MocSPh7TJKeitWpCDB2P2CHVH6IEuPfFPvkhtNkZKC6t2eSzeYbDS
Q805OC6GbXJyZnDosULy8YMSFYC32IV4tOTxwo2F4SBdCmIgVfYpBZsxNwkeaw1S
o2EMvjt4Ng+QNYZzOMwwdLQZrG8vceWkqvrV21rXJ7tnkdLT9pYNX+Z6Vl3xdXT0
caIXcDk2IW2hbsRQ6oITL0NMMx/9sFy603OCpWd2FP2dkeS+6vGTRrWrUjnxe+Xd
a+Tjamul2dCuXTca8+4lp+5wyuLCx/NBFOJhjOhXjDdcZSEFau/zhRIpv1kQyNTn
FOhgG6JW4WmxsQEzKn088MqPI/GRPxqaUeC3ScqFTuRNFIm0lG67+pnaH6zBp393
tw/VOIwQA5FUD8zIPAGZJ8+8qQJtlSs8lXq0mwTk0n7I6/6u6URao+JDDVeNWzVy
3ZIKyIXAHhQIo1DLSbouYL/6FrTW0Mrq4Pi49s7L0YoYjOlhd0+VIREDN1Q7MkfL
R2INZX2zmPniPIBFIdMQi0Z5R/B71sE48Z4yWimZFTEchZjA0xSx4sadcIxdrL6M
iEVU+tndy3tWEidVm78pizffSew3/OCVS3++BMXlyUx+i0op8cL2unwCWPZ6mViy
dNKSixFrxyOTqTDtyvg3bYZJrdbtlDEq7aBLZnLktNLL78CA2eAdMdZ97lyE2TB9
4ZODROB2QQrFmsfwsadPX6bnLNuTfRW6/XEMQ3hj8U/iHcHNnQHz3cgxv1M3+dA3
x7SMTZV8A1FwD6OfH19bq8Vlozxnys7lz0g5nh/9wS31QQlGfR7C3Pv9QrVJkOaQ
US7e3hPFjlD3ZV2hpD8uMUmquUpdQBGzbAK6fAooUi15rMxwAXSIxrGZdC68ub1O
x8Jb+4e5CrutNShcdMUvynoDb1tl0CFYhomm/G6sclNAuvjzlrIk873qVqOKuQaf
nlg8v6fEpJuNRmFgYyWElpl4TrNRmBjXR7kuZwybM7McrfY/AyoDvV/yvznTMJDF
UXfKuPC+HOAIqNfNEzJCW2KGc26Cl55j1fHmMgMnUSSulXh+Io426eaJeufubLfq
puoN7kUnBvO4gTLMrCPWjssz+jBeAyOg9PSZeB0a8zKObus55MZHGhBmcb+OgYts
w8dRAZ18V7Ihre5/Y/qwWf4clVlZUqHZzfnORq3/9/1o0JtvmwLe4PTVxBlAbkY8
O0CTgOyfOFyOxkcRMpd8oXsfHRI7Z2T5lSRP6pc1ixspUKpaeESNYzrwiwfyFqM8
gHMPRwOp4IFl/hKI1dqqM7LRi82vyd+VR7Ti7PuiI9JyZkcpzNh5WLSTuK8cpNxC
EhEzi1rwP+rr/JUcqE6DhaZCywOvQpGUgZDq7VxDKzUEsEDmnbBuV1IAJj8G9xNG
DoIy+fX35saFrR/Oetz0jpiV7fXKXFMV3rKv6bh1TwXuG7bqto4WNMRoT/9mwf6y
fEOklUcSOFtPUchKQvSwgd/ewMSWXGfrsdUuEQ0ddU7yOI6kGubThAfS0XJpkUYe
6GZk7DQFfE7k370vFMQwTr4iDBgYZHLP6Cs9qQBzlDV+1nxCfuM2uCaw5zyyA2a2
K+LK+LgOTWLV/xNQnB6J+fCgrG67sSur0PozqO/n9wj+IUR2MYo+RzRy1OFHl2L3
bGyjcDwqt+vD5t2LqcvY0gqND3DyUAVjtvGBpx+80PKdsDnv57H1lDjNZvKzHNVm
SPSDCCkJurP7tG/K394cE7y1ZP5i4BQ71QpxRQ1BGNrE3uDU4BxIIuZ/77v9hUi0
RBJtLH1RWEP2I7D+IaeNq/8JYU+4986ISzdysW+aJNobqHLuB+djKSiZqrHgq7tD
jRmSNXByBSemiIpIlYcMUpXx2gXjCeKPBhfiNb5GaKblQdP3tTvKFAo0hf4xBHgN
RpdmAWasEzyo+bOlqXOCxpF7ji7tpSQDS05k27r02j9LISVWGI1q5vjI7ktLWb98
6WKppaJA+KiYYPnvXwGTsYFwGyaoLK5I9XGD+7Yv/f+cT2/KpyNzd18mXVJXckXE
sdfIelp1sIHK9yzfIcj6NNZpgNcTChicopB0A6E/mH5dGeECdApeZHdW98pAV4TK
FVq+/LVcS3ymWPvun8QdpNPEKsehsCwnyIskpMG39cqrD7ktgTw4vwOBgDn+inpU
K/W4b0NbQbiTm/LKOCdLIG8WzROM8ZKUykYFOg4IrXKg66kaCJTU/ER8zYbA3FdO
lB9l972TlSoRrCSwrS5rEjroVhTiGOZvyfWeCuQ+W3oDjN1QVbpXPlsGLJOTZ1Zc
9Fx7L3pX7zWpnuF0eKpj0PuE/6fnyqpVmnuN8NZ8CFR/DhT1TwtJSim/Lun9+eaq
Qwm5uIlhvL8lWBCGMTbeQOCcWbCCWDFjAN1auuJhoyPgT1B9V8VBh2mlGUuc3l0+
huPFAF5xRfi3cnwc89GHwJ0JOqo2FN6qzUPutoqbeD6aYmDYeyOmEioprIuCe/Qb
LAETq+pLSs+d3cW66CW2ENwDGwoJTuTgGhykrd7vuRKXzjZo+ye8vSwMhZ3albam
LAvLCg4+UJkBr1gWGENHkk5MndB1lXAJC25NaoL9YpDHBk7+wQTB7VRk9jK8d4xd
mdsB46iXHMvKjN5N2LybFaCKwc2LpBhYuLa9iqOnyp34F6adv//l4sHHMt+jVQnS
+U/DBCtbfh+NyKKfCYmIN7NbaZdnLKLSF6mMzc9krlFOIBRiDM6hsdwmqFqGl9eP
1YnLSZd0CC3c35YdOy33v9DLjOKbdyCQKvYo9s+KMIajmAJ/BmiPnKCD4p0dy3mM
RCRqzJGSKYm6hknEfQQ/8ms5iJZKL7MxBgjk3nQVHEnbZp0lcVC+kypXBtDsNbVD
uth5Y4GVFQHaxDqcUZ2xzHp3DWE3iNBXWkh2BP6cuTJEdN+NGp8pAOuE8BH6zFJZ
XncddADmj9FvWlIaysGL5o0WPZA5yq69+iCS1UpJIxZRip3Vgxg8j3uLNfKoCGHT
6efv/a61hDqLNhNpeeBfv6oM6JrRP1d9XxZL7/Bi959NE9ZO7kcvgsyPNO4Wu9c9
i/AaF0xtbuaG87WXWSpsd4qTyGKikRPNV1tu0btvUQX+EQE4Tp0NP08mNuys2WCY
Mvr9XPEguGPoQnih3iKH149TIoD6ItKliX4spRCnRhIPsBkubiDOhRFkzmXs6495
BqfQi61xGe3eXJY1PJvULdIACGCJxJ5HTk5InBdWTItcCAb514WYTyDaqrtQaQgw
HkPI7iq+7L92Iy7dby00tgR84J+1VUfTjb9Db+5rJkFSQ2RMTE8rV7G1ovRh6DhW
x55Xi0PuCKi6plLyUzhQ0wgNG2lGWdYmFSaU7wOw2tD0SchOxG3iDbp2JBl6WNFW
ml1Y+jwz6zlK9lVNLTaFDOtga1E/xb6vWjNKVFiLf9PPjwj6thfccdcXH3OQFyd1
YOgyYLQqbA4j2bV5DL+B8YMGeg9rdBfux9vC0TrI/kBgX6uS2jasc3njNCqdVZLw
2KBkHIRd0QypW3G0PVE8tqLQrasSDV6E65NpOPT6j6/DFTUqOeLpNBuulpbIN2Eo
RJtoC/85KvgBVbqUAzL3aLyo+MSRVh517/chc6w9B0b/wDG/l3AmTlPkoYDe73BG
dR/Yvi8BFNSFCFfPEIm+pf3SY3gsKhRric0Ds5G5zG6CFubNDZAqPnNut0lH1SaI
5NSIiWek4VrK+F88awIKFGd/Jpn2STjkbsXDVT+AdMnqQQYccuJtyF5wH27yp+Te
GgTpr4xJQrqLYce7sLewWjLVnWrCrTaWhqSncW0H5aT4+7X0A+ZdkXPRNp8awsiQ
SQjwH+Gghhs10WpNU/KEOjeVuBPSkRxltYtSGe7fDLnm4VVe4v6r3TAjQShCAxIQ
2SIEPk4pf3app7TiqEZ/5qzkAuTJ05JhKvLA/Ag/iHuZxJ7hAM4uol7qQDRLp4ud
h56JQv5Jq+d2vL+VxJF8wcTOmAMwNqmvXCsVgKsu0GDP/283CdrLczOUJvtWn+lj
2Krh/9wcQ9n5uZDLRyMj99s0HGA9fEZgT2AhPXPVm0S7NVeZ5ngdUIveLRdQBKwM
1CfTIZZP85vz3qPVCJfmr6/3todsrWuwlagN1MkCTHQyBVAxNZE1Auev8qhvRdBt
uLsfwOOGjGM2jfNfTd04dpSgD2r1XvtczV6ZBaOl+RAg6NKrfLOOp4sdxvtvgyFM
VsQQLEosNHpA9oPdtlVUh0o86Uh93BCFwOrZxNKtndU3AR87142gSmnAihRHu4S3
td/nKoC64w03SiVseagqXlF6hwghKGExN+5w5sTeFNos01D22IW09R8h4k+616yN
1bGqjGcIy8W88iJUeNOlQkF6jAod8uDteSuCZ00noqyjq+DOnJbduFHr44n2WbD7
CXjpKMoiD+wAQEE90xuoDvyeE3ztrOHVj5CpRlMD2FCrbc4zvoto0EwMSdY/Xtc0
GnPNZLca/KuZ/ZPgd+OctbaJ/CmD9j0kqBFFhRGFsCyyUMDkLPU0UzezKwkS19aw
iC8g4k+cNq51BlL3q0zxxGZC2cCTAx5LHD/srg0gYw69FuDRJKLRcB/DRXecMAr3
TAwAFJ+m8BeufYh3cTilHvRWBNVxFSUs7md4JhBndWKrIL4Jg0gqw+pfi7EzWM8T
eTpSijZUm/aB9TL+U1phIZI4Tuvf8gbw5NTg1Z01CyR51vqhwt05XT20JcvBrbQ0
PTbT9N6HgKAT8P/wrYcXXMp0Nf3TiKFV389wG9fpIyemEoUqn9r0/IWRc3z/3yJq
7uVWWOsVss/3JxEMF/r7pTLweNOgOu0sjJfrp2HrrkJPx6PKztlHblBrjKac58AE
vhOMuiiPXV+5EtoU7dNtlkd/042B9pJSpRtQK8kT6c9h4r4RhMUOPPTsUDdXQPRt
015tzDedV5vK3Mgs2pRSlacLWJZUeUMY2zdwGLjh2NU40qkPU+U/vw4jvIymN0HL
ZM6hiGniNtuDtszsrOjSYbEEynKrSW0mPmoa8GAhkyszwiHjx0qv1Y5kgG5c52pE
8ThK/61bQul4/WmoWeMtJe3g9RXacBEihDPKLgiXvmNXFe59esihpLx+PrUyaRb6
+pNm9iLRiKtFnydTJUO7j9oYS4pSY8qH5WJxX+DSO8rMEHM5cUpyzYO1KggsOXrL
zVsLpBq8Qv1LM2VsohWHwX6p/55x3sMyDrVdIdmczPQfS3wL+6dPc7/jV3Wd9LU9
/D9rlbq8SO92/P8COhZfiKTa/+rOMdX2GUQAXiiJq+aYFIhAsGM1zKJ9AK4lCXg4
3hYi+3S9YrNaCRKOwTsG0e6Z8yirGTcF4gS+sBoF8OGDxZKUgZM7gatmJLaavKsW
yk1MPbow0Jyv82vaDkzs1At0WKWthscX2CqiEBp6Z1IZHm7WPoY0GVfdG49mou6B
PnsbNtSOY+3+OHtpvF7yNT9Gny4Fmre8qHctu1Humuinc5J6B8thmPzODjsBk9i5
lN22kgAItQjxbo2W5wNgkp1HMSpLaa7+w8zaaBg3CnsBYIDW8pDmGTaICsojuPXl
MJdwA8VmQvTIbKfcvda48v9CyO28NPw9j5sjhDVM1fbN8VKU8nYDKxKnPw9y563/
DM7BgHFaO/bsQu2x3dGtageu2R89KpqwsDcPdRamJGQVEf4+E5RUvfJf9Ie6QNLw
MGZO+qyivyFIDPnfamaLmVQOH6YqjmyPe8EJzL7710acTXt/CxjPxO+1UrI/sNKw
EOVmEnHCYMRcIohoBQhU3xWnD+pH87J8GbwNQWbHDvZMI9mgU4pEJygPFHc4sHRA
zZtdUWe7y8jW7ozmp2vzYcVYzB6IIF7PBfQ9qoyqh2XIKQrhKlFgdiAm2KLJv5uS
PB88clyQ9A0NLoKH/oGkZrH+qOvYKac/8CrjxTaLJkWChbNwbPlbQMxFB1bLm8Ow
Z7hST4v29meeVs7cYb4w6FqXzjScP1D/Yk5C75UUclaR+e5KbTm7kLHviWYBMPlk
tUu2kuejTbDIL3+UirUUy+/SUmI7c+ogcL1mzKckQNIhTJpZO4JHwzJOVTbIYVvv
aJJm96+CSOIQa9dCSEUN0V52RO+QQ4ckwdGngXeGQh08czhVf1uJHQd3Sn16zNM+
KMoc0ZLX0TxmgrDXx6HM3UsaY5a+1DRue1S/CvYQEMdaA1BwtDjLezMixkZan1tU
zp/jW89pjVTaM1a/yXn+YLZaVUIUgVdpacrUlwu8IDE/Z2or7i/qGBFfkaQGsY53
Jx1+wepAzSdOHUUOk60lRgYPGOS1aya3/U2MwLORxtz+PgbNingGnMPEyUApTyym
wXOthdu/gWGvUKZrcn7L00RD+HEZTrNFyavBHkM44boo72wi8O+KIlXY+sd7RAwb
6UnjW7Vl2sfiD/hr06IhDywQsAk3cmnZbRY50yjclM9Is/aEG5BI3BSk1vvCOP5C
cyX0nBn4R3LisJchuolTPv7e09CcLM3Yx7tSNN0ZBjasO1hJ+cTrfqRdjVokGTfs
22mVxzFKpAg02Pb/pgqz5pMCLy0oedtEjWHsmQjWMFps2xqk1GIgP06opnHAWGs5
WO++AtvfbO3BolKKTAJErrvMZd8OgUQr3BSQE/4F1uKeHLSOFbZA1Qc1R5nn9E0E
p2LAQAlzBkYMYm+anvWNou188dzcdrb5BwhJyObh0NnZPAnor2q7N45QRDtQIbBZ
S0AAnJLyJEaNuYOa1FTYRavT3qXsPN9GZuESWtTjqEA8RvwguqJM5LtgoJKwBa5u
LIkNS9EKoMbEnjSaYIZBJyKaTodeopNIp3KuUZs3HO2puvQ3W2JAfiFz907XoWef
aOTnHyOlmvEXVEikyX9+bzv5MDlEFKllUx85EIsLgTe1Zi2Ar7i+XumGq+gVPOkt
ovDszbcL+tPfi8MaRrsx7FRnJw0bJ+xYQPKvcR/pWCf/9+3DwO347UkanFyHskYQ
RVSK63SAnYeVGSSDHGHhRtzGKRa7+q1CqibOd/oa9xrQV6BzMDcQzxGrO7MkyRz8
uKfZRlNrzJcv+duDbyXAAdjG34+2Bsd8VGGuSdRgUsVUJX2pY40IS3HgcDePicQG
95U6W/GlqKvt5/ftSqFLszN7kBRBqkUDztL8es1aD3B/6ZMEF5jg+m2cLSmFgiVt
wd9aYrD3lHI4p/dsS7tJSZJ012o35BCal7URa8hiXB47YLJx2FDjWdkyiEA7aBO2
D6vKni6fXi/DJligMKnavsOU9p/AALcNUBGMERmf+As1fVSGsD+JgtisTMz2CoHu
fr6KGETcD0u/Xt0lsxX25ueE1NlpCJSFxaMTCrhcTwPY9p+lGTfPx66PC/5gjke0
a9BU3QpiHHPS8fKxgxVBHhp9yUqYAoSBJjwhKLmzF7yRRgQ+G4IQwUOjFg+oUuzW
CVMUbAhXmY03WgAB2JcMe6eG8QelXa1XOVMQ9XqLTDJGT02dQHGOXKrL9X+0kPOF
cBAtSa6RNyDpBBTIE6tC3VtO/mrbefDVgKX7fM3PxWDIZkAsk2rVZXrXvxFBd87Z
/RU92H5MT4oVjWGxGlVtmgGKklNbeg1F+VTQXFZmWftb8r5LBk3SRBflPz5lp8gV
5GRPmkS/tz86ziupt7DXT/GDEy6xDF1GODUK9Y/oxylArN+ArGfGylDSuvQp1SSB
mhMgZhAgtAY9Kaxx5Ybm/duD+pLp0U2omJC6lhubsSXfCfw4QYiNmrtPQ7Yu4QGZ
G/N4FIkLBHtUod+LSdg6Lv5Vw6WsYhVgjdPXFkqLPq2PAJi0+BLBbY8zJkneKf+h
g2muyhv63O1UWGbENaJ5iowkRVH8+FhJRqw1RHvvKuZI2fRMAvHp3nrkK9xv/63P
a26xD67Q1pT36zfkq1/DgS7X3gu5OnC0BqOMIiOMhyjQ5ilRffZY94mTL87zfMbl
nx3o9nbBpOG+9ES0efYRmDse7uuWEf44gkXPoLC7+p6um7lPXIEYVgaCihfgX6Q8
gc75Dk7IpUmBgpq+3EvWoy3COzPvxW3jZy5uXlJqWAUeQmzKrtv930w+BvgHEGSC
ZyQL6UdvkUa11MJJVaYexKKvb5wdU2pUE/TYv/8f09G5hFt14SXY/IemlITKH38H
IjkcpDjIhUrDcazMF4l6ETX9qzTyTVHV0qrEQ3Znp494DsQj0KEDzfFos+cJjZZS
f0wP7JrA3jFaZfuyqR7FpFxY6QsqdwjRdRbrQX59JNImjMJWqfI+wI3AHZSVAtbY
O8qIwBtvqlBru1VTrrv5r5wpaWkVFOvhrY7ErFWiQ4mVMsFkPMGtPHyZgiic5XvP
ilnfwdXvKPBlElg+6+5h+Cq2zCS0TYbG/dgl/t3NAOhr9HjGvcdnj1748qmGNuuy
yUfeenfBGPvasiLw/BvCT4vk3uPrbTRbYDdOe9XLzO2EEwk2TJhuCyTzTHjMRYm2
4TEQwKDqZzvATYxIJtvu4IUWhkd74Dvcjmg8N/bYQ8NMfB0aL30QUzcZXJnTHgCW
RTKhBAngqoruF1Qp59DQnX2QMy/p16MJKYXWkqHSFVBLhd/no1+/HlBZrNs4edJh
UFsn9L6kuHKV+mLeGfdTTdl22IMluEWGVwU2yP0doeu+2b3jzqD0kqDn/u6tG8zc
7qTnE2WvTixdXVXqQB/a97Wz8EEyNVEs75lxYF4SoyXqMB+E6SAlQDzMwyG0sXck
FMkxwGKCRognNNqRC3hmsFQHijWnQzJ6KKEbcNhnfEWc328Pt99LxAzgrxnP6CNe
xxmYVz6XGchmA5OmlSpvEVWyU+o0WGSrh5clhoA5yTbbrmpb1cW7GXSztZv4NAS5
8BmjGf3N0v+diSfPmQiCnh7huWeV+7IZlM6/7sBstJbCPMKwQk9h6HHX2hi8z5Fi
mY9wgch5drxkeG258uISTg3IiPNd4h+zC4dGe3nj0dg5hQpD3DQeeN0cPaGSJLk4
PK9oDVaC5Phh6DF6Xwwph5cwAQuVa36tvabtft1GitmnuWTty7WNfEy9MoQ7fS3C
G5kUMgwngoznTyT6iqJZOVqq4DGlqQYr6TYJNySSYRQKfkjRTXkZ8GXhyVhLfB1I
JON77ZrF+zQsPL4XL9pi5EdAGP2yjsp54fdTh4szQ5BSM6naxKZVSZ+/BFZ2VEla
BM7iYLuViZWeUIYrGn2h4WNyFnPSfA2Dn0ZQ671YVGqN5589gEad6mSlx8XsT71e
oOrHW3kXfidg+tjs4fzZHjquEixJL+DebR0t9s4ZhrdvjN76mc/iC3ZlrrCL6glF
92oUylr+FzhEmk9NpSziCFTcvM/I32A4mbWzQL190UUmHI23SgEHs3LzTvaE0BcQ
gT6Q7l83qV9TL7twyPPJMPmM+VrKAKnY2s01bXE+76ELd3oHKl7HNMkrqgtXdIWP
fNSbFGi0Er5pXGc2SwpctxJd3rmFi3IPnjYFS3SQZrhKM8z5Dohiu24oo6ghbG1j
Vk6wyNvXU6uiL87/GAyYzPKfPHbw4W7N0tAXZ4ZA8ckWsLIOJjdkNlvi9tUIe3yX
bCU9tt3BeT0nYntJceY9tqBgK9X8OWCwyCzL4VAxKbpYiTqpbwnfZUsWpu1zh2OQ
PRcCnq7oRO51OwjSqLzQiLvhq4djBOv0MitQLe9kJGT8w7E49L0jBKJafGsSIHhw
F0x4GGuOl6NEqubk7OpGSj/PoYU3q7GXdvWCgq7E/eJLcNUBtcM1wfvsng8YxxHo
O42y/VjgCgYOvjaNkG4ZkaG5kRp9o2skVFr9kdVuj7wjSgaldkJXw6FxSARJckV3
l0knsgi3CDnqMTXfCV3tlaEo3ktJjwTrEZR04A2c0ubw03DBshFRNPD27FtCCgL5
D8TDGv1JDKIteVjmr3v6L8IODhjmC3YpIYSuBq+FUdzQTBOkvEAwDID93nOoH/89
DWXUkcL2DV6P6UDkFWLXSPKvP+DtrbTR9RfVezLBg9OhmfPSzw8sBTR+EU9P4rmq
IzDQIL9OKbL12itdd38iM1WvnI2gEkHkEpP6BSX7uwD5EZT83UPR4N6qpmpRSsiF
r6LDxrSE6P/68dPFGo8EVat0Xvf0CnaBny9/aUT8IxObqfo7GcSMWdlh30mUJkkp
e9Qf/Uh4aFJpliWREg1y0Ui9EL2Bh77mxVmdlz/eixqLX/02VhdR8Hw4YCdUrnIv
ztjabm9WlJRcMrcDPyPlXUzM+OzxBGI0sidKeUJ0JWCwn4BHaamesYekAlJ//l31
jCIIl6goOwFfiMmKkd8IwPIZDYeQP+CXhpzCl9He7Gxh9ko0CW40pz/VNZIugZdb
OTKGXt9/TF96T0PzJ0U81Mo7ABvPdAfseeMgyQ/OkokT+3W9I0iZ5638yaRpGwNH
0pJRWpBDWkRlynZYifKpgzov7ndqf3yWn7hXqCPJQwH09/9dmMGStOC9HqSJfBRZ
JBqtK42bLwLAxwRmLePiOMyQWdod6YxIqf7q5ZJ/V15m9lUheNSVPmfrfruUJbWO
VNmSWAERDcyRkHjNAqHshUzEqaTYyTWRpM2ZIc2XrD9nIs/r7VpI/bVJZ8HxRO2w
mGvF1hNTp+4I3b//RW6OQozKf68+Nb/njzG+gWmgo17rtzJffhT1Pla97MvNP9HG
HVcLHpdJ+dEs8RHFhfLWcV0p4etLaJNtxEJC4PvMrt8/rfGItpFXJgP9NzFS3EfA
rL7NwBaXp3FG66Rf9rQrwpRRjh2UuU8RsDam6uO+ERx7QQCvkqIqCIO7zquqw1sR
fjDJt2i/EpAgwZfkb55lBrvkWyfLOeYayAjpZ47+dSCpcwnj7NGjYZ5tXVR6nC73
4TbSte/9O8bqmfdLJeFgdz44aqhiEnGHYRTgZTrDw9+DDPSHKn+YqTIOeLVnPHXr
wzvoz13gsAnAFw6HRY50Tfaying6/OTSuBKVr+exzZALBWGTltiaTER9l7vk0uZX
leC0kREfR+rlzqHB1gSaSk+Pqy6oCKP/ow8gK9LaLYIC5l1K74+ld7kBp8RMwkZP
2auFKOQlpW+s49PLe4RuUtmLTmmoY/PSPAK+yEmOGX4hCoiACDWdW79BAh6Otg/s
NwDbQtgkfrA53nobNgaMZjaGOQTYb6xqI1pK2jtA09i/Th5l3Uw4bfAaGnXOScxB
oVfggM7OQOqJUjeqMmACLhkODNihXTCg+Cfb8cBv41no/ZpcPKfJWhrNDAKNWupR
LfLXQjCbYjinY67hQZvJ/wJfT7x82gykvFWdiF1enPH1AACrdUChc4Hu9cfVOCXl
NfhXUBOtl28fvMvOP0w5PNEeatjg9Gp5ONiltspEGbAobC2f8dqtPMUoHjX1bS7O
a43Fgg+ulReS0ruLUggHuixlhmJrNPc2DGPrSqaN+3KnYZ2fnityrtdsAF+ZUNB7
9axayBmDK63YNF9K+MoLhGC7PHCwUEe1fUoWa/hfwdn21JV1+xcmjM0aZScjyLLq
yHTX/gTKBYKf56cU/++cxbOnEeW86It3DNFf4SeG4TNL6b5Q+4j0IHQ7R3d/YmIZ
7WB5nTGtyXagbXAbJLYqG8yEwXAgFIE1uZAQjOkIJ1prWFM9at8x8E23RB168bR8
1bV/4vVmyotuQbAxlhvR8OstsFsB0C1L3K3z3deHTazQMmC4w9QnukXGFnCMsYgQ
uusupbGlG+v4KZvTGf+8i5dO6B8zSbInZ7Qo6TrWA1mvwuBU4zRn2vuhEekHiXXM
hpMs1dZRy+Xy8BRvS1CzNcC5X0nBRJbJS8HDw/OrJ3U++3hOKxkZP/v7lphVZwco
g5OE5tTdYMWqq7q53t7omsABZcDwIQJST5mr0cdQYO6GXY6W8981CknqWb+DwX+T
wTNP3fTdmc+HfLYDXqKeTWoJPx1LlyIytRvNC4AOPpM/xM7mR/tgAn31qB3bKJi7
09NAcxW9bhoyILyIY/qCApnOx6ml7cXL2hiVCOr0DSy1AJas4r31GGYKZEzk8n6e
fNW56S23PewzNdr/sEia9D0r+IvEDzNzExpc6W7f0E/cOBKCkThevaA6tO438hbU
FiMg4O9SJASbg4039Ekdp3DJ6Ab+chI1/IKxKoyTaEA0G9gMh/8F2eg7mqJ6CS54
FqSSJNtya9eckzVKvvWzdoXUpUe8q6O30gi/VhQrAhBEX9c6QbhLKwnu5lJVzzb3
1H6s5zyswITM78gs6hxn2ST7z5V7QtFjvB4fyBqOXtitVK+ekRH56il7xpa3g/w7
4vVV0k9Yi91SwZilwiMxMwMGCWB139S6OgIWXnDm9MjyeofFvqJexj1EDDDkLgoe
bPmlsCh3MpbkrP6r/zcbSRHTtbsO6h7YEwaJFTK1fQQK/8MHKbvmGko2UOjU0Kae
4IuGsUKaBunbG3ukIG5inikZ1ZijxPJYHV0wYzFxRFlWq+2iFxnjknkGF/ouBx20
Qrd9Zz2oyvkw5kIatsmvqwIN685DiQdJbu6Mp4RBZ7+1ZBszcrmDXZuVj2MYCLnw
`pragma protect end_protected

//pragma protect end
`timescale 1 ns / 1 ps
module `IP_MODULE_NAME(efx_csi2_rx_top) #(
    parameter HS_DATA_WIDTH = 16,
    parameter tINIT_NS = 100000,
	parameter CLOCK_FREQ_MHZ = 100,
    parameter NUM_DATA_LANE = 4,
    parameter PACK_TYPE = 4'b1111,
    parameter AREGISTER = 8,
    parameter ENABLE_VCX = 0,
	parameter FRAME_MODE = "GENERIC",    
    parameter ASYNC_STAGE = 2,
    parameter PIXEL_FIFO_DEPTH = 2048  
)(
    input logic           reset_n,
    input logic           clk,				
    input logic           reset_byte_HS_n,
    input logic           clk_byte_HS,
    input logic           reset_pixel_n,
    input logic           clk_pixel,
    input   logic                       RxUlpsClkNot,
    input   logic                       RxUlpsActiveClkNot,
    input   logic [NUM_DATA_LANE-1:0]   RxClkEsc,      
    input   logic [NUM_DATA_LANE-1:0]   RxErrEsc,
    input   logic [NUM_DATA_LANE-1:0]   RxErrControl,
    input   logic [NUM_DATA_LANE-1:0]   RxErrSotSyncHS,
    input   logic [NUM_DATA_LANE-1:0]   RxUlpsEsc,
    input   logic [NUM_DATA_LANE-1:0]   RxUlpsActiveNot,
    input   logic [NUM_DATA_LANE-1:0]   RxSkewCalHS,
    input   logic [NUM_DATA_LANE-1:0]   RxStopState,
    input   logic [NUM_DATA_LANE-1:0]   RxSyncHS,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS0,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS1,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS2,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS3,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS4,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS5,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS6,
    input   logic [HS_DATA_WIDTH-1:0]   RxDataHS7,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS0,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS1,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS2,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS3,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS4,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS5,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS6,
    input   logic [HS_DATA_WIDTH/8-1:0] RxValidHS7,
    input                 axi_clk,
    input                 axi_reset_n,
    input          [5:0]  axi_awaddr,
    input                 axi_awvalid,
    output logic          axi_awready,
    input          [31:0] axi_wdata,
    input                 axi_wvalid,
    output logic          axi_wready,
    output logic          axi_bvalid,
    input                 axi_bready,
    input          [5:0]  axi_araddr,
    input                 axi_arvalid,
    output logic          axi_arready,
    output logic   [31:0] axi_rdata,
    output logic          axi_rvalid,
    input                 axi_rready,
    output logic          hsync_vc0,
    output logic          hsync_vc1,
    output logic          hsync_vc2,
    output logic          hsync_vc3,
    output logic          vsync_vc0,
    output logic          vsync_vc1,
    output logic          vsync_vc2,
    output logic          vsync_vc3,
    output logic          hsync_vc4,
    output logic          hsync_vc5,
    output logic          hsync_vc6,
    output logic          hsync_vc7,
    output logic          hsync_vc8,
    output logic          hsync_vc9,
    output logic          hsync_vc10,
    output logic          hsync_vc11,
    output logic          hsync_vc12,
    output logic          hsync_vc13,
    output logic          hsync_vc14,
    output logic          hsync_vc15,
    output logic          vsync_vc4,
    output logic          vsync_vc5,
    output logic          vsync_vc6,
    output logic          vsync_vc7,
    output logic          vsync_vc8,
    output logic          vsync_vc9,
    output logic          vsync_vc10,
    output logic          vsync_vc11,
    output logic          vsync_vc12,
    output logic          vsync_vc13,
    output logic          vsync_vc14,
    output logic          vsync_vc15,
    output logic [1:0]    vc,
    output logic [1:0]    vcx,
    output logic [15:0]   word_count,
    output logic [15:0]   shortpkt_data_field,
    output logic [5:0]    datatype,
    output logic [3:0]    pixel_per_clk,
    output logic [63:0]   pixel_data,
    output logic          pixel_data_valid,
    output logic          irq
);
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
GSd1xavSXoxmRINmTKZ6r3Y6Zp0e5DPK/J9d7CI+WZ4BF8cpjGIJKdJ+8xfH99Ta
pD/b8JNKD0mSXrvg9Yzjg9iia82goTX88bPCtHJqcMWxqjYCZoOn/D1yOoHL57Sm
fp9ZSFPzFb/mdDJvZXfJsxaEXobv9k/4IKk+OvPU+kA6ktkM4RNqB1KCTcZRFuQV
bYQ/BwitBJQplGAJcYEUJ/DsnRNzQMEu2MiDsxIxMQdyyjGHHEMDaWwhTwsZAXHp
1K/PQ/0VnLk5N/KQ9+lVDopy7Ftk0cdpH5sIoV5JcLQeg3J8rDYhsegWFYdWEPPf
gePuHCLAsNsQpQofEHFrzQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 19520 )
`pragma protect data_block
L0kUbaJthInVYQUvrq9gVf7sP0HnhdfS0KoPQTvnt0Enx237gUCnbtxr0ica/Tnc
GsIt4YEz/cqypVw3AUVd8tYhPPgx8YtBOcy5m3G7Z540hsPzYGhOdKJLumKAg0rv
0bKtrUki43YEhgb23ekKOVD36H8Rd1ljFuxf17LCRk8nTljlqjYCNFukKXANPLA1
p51TedUgJq+B3xPWH/Dhcuj6y7tH/b2JnpHdunKwxSQQvEtsLfZaeFh/r5aV+uvh
PRjjHUjjpcceckUTDAPX0bRsZ7X52JvJXnMxJI7B+OEoFktNa5zKzzQthUUzLd18
21f1zakAVxLbGmPH5pUzxTn/jMKa9Z1OQmazk1xKHpDQMW7PAI+/JzT3yXpHcDr0
eygndWKOn/c9KntHAQk7Sxn5LDjz1i40F5CApqHVQGIoHHxBV8RJrPDuP11PlI/x
OZRY/7SA6WsmqUqmZVuctjbQi/QhnX9bQMOlyN6+neJxZ3XTNJmrxYXNbrFey6oH
YZD42MydCi1sh45s3Lf2d5oJuwD8vs+e8FzC9lD5dMPmJfjtm1Y9vKpdKvH7X4XD
UzcnhwxMFZJp/52p4CxWE9d0q08ZxvoW7S5/fGJcSn8bccqyezAESosOSZOfb0A2
7N2mOwzMaBVYEL4tDXwQCzHhtCklJwUiCFgXgWfI2016A6rpV0hOse4eT7pDLaEi
75ZUUE01RSdZ0halxSidiUj9v0Os7aJUTE2IhQDihOacWk0iitzP6VmWkTevBzIZ
IrkkkpNwvZE9pbIhbMA5fx1RGOaiajbUkLIs8B7phtsZpq8EAsUa/BDAsHmpC207
r5YPwq1qmgGM3FFDRDYS2EA7o3ALgYj/1qfu79bjcDvV1WwKFZIsFQrA0gHQ71fS
SZcdJtAUEwbH4XNsSi3k5s6mxnrnWSvDs7rEFrCPYSiU1jW4eKL5LYM2tYdzce7T
XHDymnA8Ktj6KvHEpC1Op/u9xOTLWEVLQFJ9w57qVsXAhQifa3CnqQwCTKBYSgsh
YD72IfcI+k1B2OmO6MIWf+798PP6qhKO0tA3dOTOuUqEDnQTsnfiG0034s9EgGiV
PZ2hVUhQfc4gUhKp11q390ie/gmgSBitzQ6993p+J+zTR/zlMkwwTHKqeuPMp8Nx
T2y+Z5/SQhbqnnI/Xcjz/bn6R5xf9D8m5QZLgnuL34zFaXXPXKcHTdWwO3Ii1fot
1F+bQAaY2ic3mIgt0aAggkU1U2aZSIgDLJBd8alzuCRv2mEuCAweQx9FlZBXdwx+
vHmUKKIoU6am7YsOx86GkBKwpB8SAZjag7ir8Wp1PdaOvuVdSE5xMopCXzcibMqt
G4t6VX9MpgjLzyv6U4/mC2wHifxLxTd67HRVZGv+yhpFh11tINxbGCMEdmybD244
XVJX4/BIG58LBL1natGFKJipX5/xtAPZ14DSSa/oqCyKd+4zmii/lFROw+6SLFSm
oa2+cIi/xEiGzu226FV8YQH2Ce3P2gQq52f0DyMiJHOCPHdqsgsOmV9IL4Ptea1t
PqCdOP1xwqjLZjqlL7ayYw/RjfeSpMrLqWmgLYvYgPgG35J99uxcI1Dmj1wvfEzI
xJVWSP96HskfVFogGQt7PTzoFBRj/btwnnauPkRIQmZqgtPTrKn3GgjmHcanhMIe
yvIGVMz1rluVjgLMohrA89bX7Wj6rW1UZOLEyXs207QeDfCOHi81rZcxulkGQkJe
unPCZbezgPqYMDvLBuLf/lz4UZ0IBLuoU4SC7McQ6daq1WbGT0S5Hp21aLKccd5l
QD8a/ac+8ZOcYBOEN8o1Hf6qAXrkSf9//M0zXz1a+r+SOrUx2VIJgxMZDX1EfEat
M0ka0POhoJHYFagKm6dtXVnZmG+0vWyyTeOiAnyBILFfZdf8YOYjcBf28hrygbxW
Bue+oybUytCyvEixTeZNVE+rvHWv8FeSGRIk7b1a/QI0R16kLBp7ZK/XMLHH/A/O
H+INXDHAXji5pyIC7eYNpbsVUkJ9uEP6YPTXSl5V1gq9G7EiLOvD04iB0IxjIQkV
AH6jL4mvVRi/Fk1N6eXQZEFVP2ZUhlS9iefC8Vvsa1xtxJCOk/4w9aQIC17b8lyc
beOoUCuuUSLpdswf1YuksGTaehEsUTOOSppz4e491DgAelHRRB7gKHl1AqLVkJYK
TReo1yR7VKSCZ7fqJigXbxhB+a0qJGyIMHmoNL4wkA+muNlA59z7KF6YbD7ujdTO
hNrC5pHOEnr+y6WLeYe4dl8ZjX8nxtiuNt2WRqGGyrBQocFtuIf1Z90LOrw67RW8
g+U8iMkBvvoofLm2ND2/ckviUzoJOFMDhgyjmokASGckpyktfKx2qcZJECug26MW
q5VvMTuywCjpxxALr7aI3V0qz6LIyFMqkedXWOdkgbTBuerKnc4jWgjAqyBebbhT
xPZ/a1r3n3mMeIP4Fj7Z2pfItDuSwgutKj/9BhEdR2kzZbswUbrH+1W4+7tbgTzq
gGm3gVgHo64MGDrh25LubGvnz/QpO56M3I9nkROk7dZ6ET3o4R92xmfDjvTVUDA0
kkdq2N907Cc2IvNmictoAsaF+tVV+ryrZvDQQislt96w66QJzCIWHo/xNfHGEyTT
PUePh4zfnHmbVvkqDjyP6EGH4keworiTbCSaZq+gEccW1z/vn+jDDijY33RUHvnM
S0dAORdXRJRnr3S7l7M4j8xbnqVhKtFTTLY3QYESqhhWSEM780ovG0Lsu1FlhM6/
t6sWOPyibgobcLclvRM5RWvJXk5Su7ZwM9RyiHrTl8wjpX8TxcxgZj08skfOQkpj
D/WOBzt2Us3iR381Q/eVdwud9SBYAAIFdNuxRXLKZ1gX/VUe89mOj6J+KJUmlkU/
ZuRJylD20UP6QnbiGOneu/JOjp6r02U6BqEXV6KwrynqyonDIF8CPWugxA4HOXzI
sNNy8bQF2Pi4tKpbVNNi1QimT9C6cbxjrhkuXQREPAiOwaEILBUcnFHM1EYXJbgp
mrsb1nW00XfoXgU03bD9C50GNgjAg+a4+F8RASMAFX/XMIrhkMbYHSAGZaGzLuwq
3wSelVQFB59BuQ/U6tBFW1H568uSPUNZMZ2tHCocc2qrLZAQ6JxYx+vWgSMqwZJd
mazfHsW0im4hSRZ6lffaSc6xApUbu7qGWypXuAWOySQlQvDQE7O4D0CUp+A+fGPy
Qqbt4zOzBlCIJQUX0EpXk6a97qisPaw4spZ8f0sbYo5JOnFjvFrmTrjNot3AhRxP
4QT/REJTe+3s4EoCDn5fdzNH4YbXQ359YSHw4TSGjhXSFDkcIb392cmKcvLoErwf
dI/xXYwpvN1ALhoiMq4475UCit0qaQmQh/kAaJwOY6BMvMkuuZd5alLMex0bbR/K
GLJZrn2K+2hB5hCSBJeMHz4QtsMcJthDSufxaRAVX7V3jFcJsp9Z83IiRl/wGOZD
8JqdnnyY7qyxoMQ/HtHP80FE1Q0Qi77I1cmiI/KIUKwKyDVSxNlhDrk0Xne8vl0l
tsUzj0TQlbe3W6OLPx6gYDPML+OWqwrsaJjL2WTDDn/5RWJOCHrkLe/gsS54OxpQ
i4It5hosYXslC9dTZtEiTWcujrvKILXxUMhWs2VV0HbuV+4LtM1ZzwD85ztnTpic
XH73TTZIOLU6TOw6ZFzvV+2yRVQyNXK+r9BGOkR45lbQgQH0yfliztxf7/dKH09D
v0Rh/8btjLo0oASNP0inD4Gl9wNQV1NYJUmuCx4H7rNA/iR1W9zbHZNfrnbQAXCj
3amPHN/9c8suAopR0qlnwQqw1CLyHok9QTXhB5Xlenk1y1cZMchPBGL+kilHQO/g
Cu0u8D7yQ3Iyj9oXL572Z4D3bGkHj9OkWSM2v6Nnysh83031E+ftIQa7iEAihWw3
PRue3tZVNXz235XuFnDe9JG9Sl3ZCMZ8KhS8juyGXR/sux9VsjP2P34bn8XiCNqP
QjDHVPswPCAKNoAdaccalQsvGdaTZEo0stAox8cZ9cPKRGWGOS+ZCoEBiY58vooC
vBn9nS7pEXds/WJTL4m1rkq9gULnSacNHxoDdZAXOI3ockoDyzprBqZ++EwcZ3nV
aqL+P+D+0BbRTJM+CEjRG5FdkjAQdb6oir7ASENMyaN0HDtnZPJsM5tn8vJOj60L
eaWib/Vnw5eS2y9K8Al8RV92OGjIAAdUX7PQdugsgHBuAE1xvtMttJnF1p1RXHMI
zJOF+fUB5tqAYo5ndm8cHyfqCx9UuOsX7w+Z/2LYqkm4m8OwLw84a5L0LCRPou04
TJgaI06vcep8OSq0m+MI/w1fB9JQ/eB1t3LtY5SKKcKt/4P/4gGjlDXHxKxa99/Q
/M7eSs42aNTbjpzI0SutDw5JDXYF5QlJUhhkZB1XErpSGpOTcYfX1BEQoFOKV/fs
YIlQoK093vnmbYHeiHoeXYfyejEUCxVsFzfjwAlVfgYXBFAlnrDHwjX8ctXb1TIC
Ok/Ib/OwEGJyUn3aQpI6LVNIVfrETCLPFyc5JE631l7xnweM28Lr+IoFRlObNBb4
1GSemiK4ZIxTwnFxnI0SUJYdNPaYg7+SgNQ0ii20edDnh1fn/nJf3M5B1VuevjUW
eHJLz+c7fXZLlb7HhuerHbW4aVQ3p+P+03G1ZfhivthwnnlTkVE0QtGzslVxLR2i
y0QbLNeHExR8HCcAyYPIKZopqF3kdsrB2eH9VSv+7D+jkmVsqP37uH4mJbyK6Uwm
1i5/wcTHu09kI/jRSOLKmJuodLUr4B77H4GBM7w/uA5Fzbi7J3CzsQ6Iekd0O7Bu
1gI0RU2PNdxrnnu4Kk4curNGztIdJFS6EkczUZnnyRrekcDwwXq2FWUkbH0HS9Lf
CkQe9J9fcRYlrVFSJAJc0A1tVbP9qv+je6zLetgEsn7Nsfo4x8RHDS+wI66y98BA
JqzXKy+eCDHwyDIeCnuxn4PwXqCeOl8NEXkVbdzuv45SrTvTDuxK8GCfgRohnf/V
fXnVJdB2DmXdncuikmGdDFspkMcXuKEUT1pMijIZnJHuhVZ6powJOAoyyHOyjeCS
J4/BIJnrcRtlnq3FfrYhS5InEmOcVzYoii7wWVDWIbdvJZvm3dKkaPdKI+JQInFQ
Kw2YQwulX7G8e7D7lzUL3Fl7C0LnsMiCe0/d4qn4JeJcvU3wHyyKnCSCwM/fjuXi
maU2VSq8NGBHXuxw0KSA1K0DoT/Z2jgfX2WaOjZRRn0PRC3HvMh5cdqwhqm8ZxGa
idfxgV5NOcLcSVYkxllJHrX8OzppzannIe/Gr5X6SyVFvRDcg+9ntig+t32Dghww
xZS99bIu3YVMb2IEP/5TfST90aPDEQ95ik0nlbZLr/K3yXgzJGgac2R9Tyu/Kuhi
ETwKDYVglGA8Y1VqnfitfcT+7C7ZyTRuq9XdJSbbCAUDBs0ZupaaUSqHAuarecQm
rrkk66lqPg/Huai18I5YR85s0LwBUcrC+1R0AqD4J5twk1MoBvdUJHCymr9TR4Qr
9hc7sUrJYshUIIZqCDPhXpQFB+/f+J3gbK625tvGLOQBxupykHVGrG7fz9m7//Yf
dqikM4jWq9zyVMuoDHjx/KTRyXPzHbFKGPDDuxDWXy9yq4rktFJQt+vkQwpTSFvv
ispZCPRQZZzP2qLCF5XrgoVKi7i/Ft3HdcoubrGLn7wu6UdT1TPgRyIsojNq9QiK
2Sh7lONeX7+8gKtmT0Xu9PSQsT77zJMY5CHhsThuue7K7nrlB8E3Q42QE7QZ4B2d
jFBiAUzaFUE3vCElTbylDs0YJ7PKajuPty5dWyq6G7FzFYVZnmZ2oIWhvyteLsw6
VlqqmrIvDYeN94hkO9mFQplHVmIN5lEbHjDAbFGwcct8y3Xm3BP8Vu+yiWJDpl+8
/CgQuS2fH+g96e+oaOXqL3+nWExLuv/QlrZOvPPqt7jleqPUsPlQFNPLGUzwYHAG
+TixAAUU6zWnPZYLrIoC5mhV8iiN4p74XbfytkD2BPYlOG+mryQERF3TeyFwpsz2
xoVnEqMU7uQ58Zz4lz8Hzrl+WU9SkO9IQXgn+DcrQDDFozl0zBH8m+BqA1gPMO9K
YU7kEo26/YiTWUigz5WyAhNUDz1aKU8PpPfGgWP4LhLbpO3DzM+x+gyZVNnfu11G
M6mDRQ6SpjGb561178e+tXyv2sh9qAF6cjn9Wj5M8fh0Nev8k5Y5GaqHZCBVXTwK
y7DiYawB6hr25Hm1tfpBl6KPQ6i9QlPXQ/NmDIZYlAo+/ydforp3P5yrYVq+kYyO
N6PNgrEn1kOoIWek3MV4PxPJ3DMlOyJ3g2S9zJgO4A4zfiTbJzNyjqa8y+mifugz
9WoLFUY3P5SFY+5E4rJ82Dkd06PqfcxDw86lz1UkziMOHbn0RKXkHxFEWk2OK+2/
Ag/vUG1CJVWCXMRrMReYhecevbhZvx6Izcq01pBu50VXYs3FYyjRR/1cYTf3wrjN
U+GjERaOL8d8iWX5hyYnHB7MXIkIVGrjCw3LAlohhcLGOasEar1Y984j3df93ALE
bUQM4Y2qoUsfKav2rgmKjiCblCsGD6qECr4X4eE4HnPvOihEb7OE6+VyH4KSONx2
OzQYPFhIIwkUBQvJFGWS2x5jzw+l2b5lYh7doVP3la5At2TJ7bveTpRA1aamf6zv
/8k3fTwNmuK7USIPQf7JfjeVGeAB45v/o9/K05vyAIVHob8d4O/OPBeTncjLfA7J
O4pEQmkK3/e3LXMsFLXGJcUdAdqsIhHLq+NzbgSFJg6eGt55U0NEpp0GgovOSBpM
fiJ2EUmQbngNubDAdsdALzHobYH+SmV6+Zpa7r1aQ9Ni2ZgC15730wWpoMDjFtrc
WxeyUprsPPFxIOzuPwTo8FieNw53SQBmiTMQnoW1lEkoINu2CPqIquFU3uT3bnhI
Aabh32F5txbOiiTDpK00WnJlkK+U3NvxYyNZDpKsOyHMN5Poiiu/PLiUch/bloRC
zJeHHw40PiuykZSSSFVZ3s7sUsbz6dm3JHzi+kFrOzMzH2+wNInQq5OQcRHJGiD5
Jc9lHDQlG0HMO+bUDkwkGpC/kaWAKkI0zZj5bv2+ukOvzpdtcNf8kJ1L3QSsDHyq
o9PBlnHDgQmIAmFJ6B8ISmzrsxWnZMxawv+0QgTFGUL8EE5V8dIa5Xd0AEVHUaKn
ekjuwGF1aXbejowzejIsXsI5UCM5+9tAr93SWpjDmrK83kto/D6PUBw3kZRu25as
yo7QAPH3b+tLJtQoE9qpxAwPDMHNb3CJ2hpKeCBdedD5TmO50E//VSOi2NKUQd9q
eRDhyjjqTwMDqzjf+4uB4K7cBksQoadv7g8vlc1xE63Gil41gUrLqiyI6zd2kLhu
1zsD6mZCzbJXyp+OZnR81ZR8C5cP0wk2/Uhm1E6ktNcS+pMedtEgI7xiCn6q/Lo7
Ipt0meavh0WZnTW29J5qmpGGH2UYwCFypBEVRyMpKbDAichoqL0Lc1HLTUC2RAvR
cbUQ4qGCwsCauyQFZRxbve2QBwHouN+smpv6iCGXm7Wc4JFXj8Cdu0Rla1//Vpbt
Ucg0CfazDH0bgUN18MzhnNBhUldAYYzksNSu9bzVPtrH9OtSV4t7ecZGKUcwaID9
vLfq5vPW1OKtl1rJ+7IGPMKv8HRZSzqFFD5HdBoLR93Or9qrM8fP3S3R0EZ3dYJS
hlVliT6dVWRSwQC3HuuA6kLZzb5VQNVZXKiuayaaTJgU5FCtYAhA5Jyi8hOSV/Cr
iyKecuqwa3ldZB5ZAIngpT9p3O2JSfQ8mmkyN0++rXqxer93q9dMDpShPWyvXnVl
E4Fy6YyBrx0rZiM/B8YFMiBzzQluKl+D6fBDN2hYvaA7UUQSdK7ySxxZdXwRJbdp
Y/HpOP5iNAt3iyAPqXy7H7/78ekkES3K82kcEA3/A886LhMTbkNAsJhMR2JZDhsf
Y9IuoAT+oivosmHygVtyXJX55CcrB0uCMIJaKFxkdLov7CEy/g9OHsBowTlplY22
AnWYLaVKvgz/B1Wto6hTj08XMR9r+a6NupDgeXVROrLjQD9DWhZQm3RETqhN27SR
UOFC96t+QoKdNxdoFJABKdnEL1NbwxrDOeSn3j7euSGcogY6f+EvPTylml3gDpRt
i54okzsDJj6iOe91iJLe4Ra0DWRT46COOEH188dQQ8dCb6O81uYB6ahACngcT3FA
Zo4Kdt3ar3Hg2AwCHGKr7Av0tVzNcsVEcCLbhTh2A6Q3njQLrrwdgxzR4tgzzLvK
IrXgzhEnmruDBIyLRqCOR3i42x8922O0zz+d2WoHYQsu00Q7vWDZHFK9+k0imwhx
HaXKapdu7kunQKgiZB4j/UWI9Fu4yxO71dama2v64Vj69lrxgcK93Lr3oUo3OdBv
7uWOePsyIrJj4TmKSRAq6RDFppC8ysEYOFmRgIfvjBinj+Kr4DvZXN6TSNan2RhU
0WeypXRJjbGae2e1ooIxfagHuS2cvb1mPxYmZE/TPQMcAiZFMWgR6U9zrP6ed+CP
n2PXBhpcVJVyEzQnovEnsta/09l5BE62ZNgHLvD+wLCN/Z8safzJfFY4if8VAMpv
IVZjQ8QREYmgeTSiAkq57ysMiy1L3Xsx1XTeCC6LRv0xSk6m6xl+7Tj9WihAthQ+
VUCZQleqpPUjceZcVzQhkrbbn+u+AGuy8C0g7uzLHZSvQD9qzWxh3ahx4W3cCUSE
GL1b39oqCMVDkP2IpUKO5K4917aoisY6uK6Xmj7hPVIBFW1vpaBU82didBNuFbT8
cirXjWBDIjRJs/w8gGKhX0n04KRqrR1sLDPqGGE+TghhzRkw36e17IRvWYoX/uxx
ws/9p8krX/yZfj7flwlCWkVp1US+m+7Ib7j2MFDqcDph/iRgzcRAcs0TFQTpKb68
TtXEK1V6hzWEe/73zOFPq8K5Z30UQ/oW56jgOWQjXy6qo7DaLrGSIQgHve08o8SV
RqCc9h0IWwxPxtYV85l1SgHGxujUKAkeu8CDVl+zKqNj5zoNWUF+PnOciqqFLtrG
bJrty5zjDfFthI+MYhgBJndWIOIP0EKm2E+3N8KifaehHv2OYD7F+CS4A+DHTBqV
FB5Kh/OyGdMvx1fuLcUazKcoPI3CtjvXdyZ0Wq98gSH6tCXDKEh4C+fXJzx6W7bf
Ad4oRWzVRkjr1gLo7kjrxSYM9CG8YDGRgnx7CkwM+/jpctFpC7kko080Fri69Wym
tPQwqRC1zI4+rmyJOwoaiXxt2w5XiocAM/4bKw10A/pSbl3pjBmHrZztjvKTp9WP
boIoPt2Rc+/wZJ0kz1fsiCbObN3XwyCdqva4rbg2gHIMNNaet0RQlpFsrUIYdbp+
lO7s0WIjNoKOdSQkd1eVkOhT3nGMZ5gU2b5tLi8DK31/favVsjn0R1LjRfVujjO3
j7bHt4JZH/KkbpZrWITHWpMLDs9LMfuNPER3p7eEyLHAymJ1eaP2x47HUXVbnrRD
xDoT10aDzIDIbDd8oqiB/TZMFg/ln2Y4ZXLapLU9O8ZpU0hAlf4db+36BMO7BP93
/S2MMQnrAtswNtFKtK9fpEfeTaVbFwYrPx1jEOUkr1ysrXlGW7+lDzTRy6kbi//3
MJ3z8Cj5sQ0LkXZJtH+CaHqsmsC8g+17Sc1rQ0dZGqphGK1RainL6uQ0H895gJ8a
nmFTNJVxQePnbcEKVm0ex+uftmKmnNEjdgro57EYmB/KoTYA5kcdrez8seOxwZO3
nhMUoJiG3Hlcj5SNo0GFHmVg+Vs5plcVUH2EJ6zLAlGrugHfU31uIVJh71k+OdJm
6QTbxla1sfZUDnJri+Dlj56FnmN2IRwaP21bBcT2BCYshP1zdJMKvnga72OIKxZp
9K0i1aVmEJi4LpvIbRmRk5aXgCsByTvY2lFbWaDpDMsEM6lv54Wb55HdpkM7fx+Q
ujFlntCOtcCOoOlignhzYkXzt7jY/vquwFjK8l81yiYnWRerDpIkeLSSHuwvXjk6
vWpfbsa0Liz+t5eI6bjc/CZpwKaj+/lxxvwkQL0yp8eywu6go7z+mpeawN96/SqT
NiJV4+8qfjK9bEAwUsNQQEez3PlTi15PtA/j4mYb44GGylad7+9zvpM5MuT47rzH
FHF73o+/nQlBHrbtDJiHRtOfKKy1dRpeycewEZAQta0RxGoSIlV2LtJhBc0nmwJZ
FZSMiv0oqj6siJut5zMIRldGfDQTvB8PFPoa1nJjtBD/FHjye1Uf2IrTqwxUpCGw
vuiNYRfD1/3RveC4V+OSncS/P+l+iJ2Y7uT1asbD5/OJbnEcqemjj7jNyZQF0Aod
asNglIYFjaRNF1IsDJJ1TI6PazkF7WIiY+HkmPKIJWJgO6/IsgmkeWzkMksUVZy0
GpdICp/2GKgVOl+Z8sEQpjxvT3KmdGd0KqgZ83q4ffjpTA+2JoVsm2rJj3MjV6jt
IjXSHT9nfW6ZU9EXfTeRPB+xix21fjtFpBSrxC1vMGmKnANxCKHpFNESatetnd02
uXKcvAGdNV6pQRKuStRzW9I3TUxsDyB+ioIBEL8DfDzjhY+9nNil18OSnhsOTH9U
Mem0vEv9RnUfjY4aoZCJQmICF1RRq+Donhgc4fKVsJ/AVynzrPZ+RJJUiEQDYorw
9wQMo3yDSbIv5ll1IJuA6LlSEORmfqVN2wy69EHsFZQB3I5mmPUx15V0BG98nNQN
G3IzozcfJEUCBEprQ5Xa4H16u56gzfjTTOCSbWr23gFkiXTdB8/b0q3Tnpt3BWUm
m4x+ZEc76tg3uNw7rwqAtmNLc5c3uW3BDB0+fHRCb9x2V8Z7s3FtFlsvEwwD8V+l
U1CgSdafCHjoIBBZqLbybyYu8TNhnz6DSUcfNogioued7LHr51kSRQruBDS8loIU
eIkXjF2k8rnFvjIjtNir535yD1ETrxp1P5ec2Gwggy4DnT/m5XCu/XQrRzprXjwV
WVn4yDk1aE0NP0dD6r0LXiTvHz+jNoqIpbezLwhJpEmnBAjRtltLDLcjHAZf94l+
nsOPbJrjJi9XT+D1xdW7WbbRFDVG8RwljdnjfCjotFvnN12ei2hMdCwCzk0dDQmy
jvkjNMNom0OGSordyxRgFk4pZ2vn+wP68YH8Z3MW9gund5uwhrRJfuiXwCI09GXW
ylTc08yI+s+toi3JITNCZwjjwkQq41dr9Invk3+NAQwtDHiKif5izDl911K/y7ov
8wsKQNvx9kLbXOd3SwcU0QakqQjvi9hAeGZH6iOY/9l59BNk7jy4aRWPxkHYmJSt
B/0868JtStbgKnvFZhu6m0j6MKS5LVK5/DmyvRO789qvP4MkQbgYx9EfPrgRsX4z
VkHA0Pfe2PbLf9mb9jxyCB617xCdDCXmfMJVLe08H3sTG6ohtiGfJi7j1gaK8phb
seELQ/CdcpCsGt2bxut/9TDwGXfEEt9k3hWltLYJ+5BM7OJGar3kMFqP231hv1st
uUgNii2HdLZXYIxKbP6BKpqdZo+5nsWuIdGAfw4o0dxKx2G8k1tRJwskbEfUds/J
s5gerAS6IRChsH0F8Ku4bQa0Fc+psiCMbNomni0vS1GxoSR7/nFg9Nw/3h1tosRc
Ludp7ZQobt3Q7pRsXNbpE5DVfBrMVGmqoP0eYo4GLTfTM/rLK/HBFyIMxVAHQFB/
EFGlD02JZL/4be0ucbSdTCBJTFDbyCltVkO1YsGh42pSnXc2jM628dwDJu3uagEB
mybquYQP8mDRs/1tTIwXD9rL3ph5KxTXxda4Rg0obwlMewX8FJV4HM1TXzzXyD0d
B5eSK4AGZqFEpzu1TKKNXtveztiMO0rBC2qRKE+diaPKS2NTdnCcqy5OOZbwrvxX
pMGacjQDeoozuObfjxE9nbSaThjmec8zidrpwx+pUzRsB3x9nwXsYHUT3ebStI+N
i+WaprMcwDNTigimXDygLzsyT6UO+F2lIybBid6ADIJaFdCBWpqCrpPTKSSeSxhi
vI/U3JHVkStKRBgQCtTM25JBAA1UpRIn+UR7a+hZJdcaaNKPufotac8X1Kt/4aZ9
u8hjepye580/KjgrBFFv5+rQtjik9VYg4lcILNWpr/xgtiFIDO4p1dngmKLFd+TF
cFqsfSQAcmhtFIiKglcjYACHvW4SZleRBAL+rDYDz9ddMpg3WJioTMkoHFuNDRpu
fbUkiJbpJ3AFpL77hHeqRBKwo/rG87nvNO/efFMPi0zUlJ4qh/PP4+YQIWCydtjk
RuAxR0rSfKs70KGITX37UCZaEuhdnC0uc7WJJ3eCSmRJuk5BfNgEKzWrp4iUNEWt
cuXVJ83HpSiiHKjfEv7BoH5IlqkA9nbYdXLunbkn837ezx7HgRmtKLBOX2KiWXxJ
HEKImgGLhMO46slMxqLsBeNx694F0WtXpOq94SO5ujNBKvfqDPXDs4mQS2MDqJMJ
6/HEXRntLG+Enry/MrU0ma1O5yltB1/+FaK+3JQvnXGrlRVuKxwWDYQu1mznQsLD
DLVNrxXkqZ4Q4tghq6ghHMyENpuPybLyIwTvcWBaXIWhNRLWSCcVlA3xxH5tVOMW
ocdGFqU4qfTjV6ifvVlU+sYWq2TKIklTEvO5TYuMgXyYFgVCU1qPV7AJFFGObqZj
ZkrV3mL01L/Pv+UmaMGUUUDWbvHuPWcZohYe0ijN0OKK5t4T35mdLsEEkPqdGxX6
uxRxrdneRVZTL6y8zVfXGB2KJmWT1ybuga5ti9OZ+qhXBeFzE4Gc8VtI0tj8InsX
WD/JQ/6qUoSOu3JPSqB0eU7+aAp27t1jng/i4tVzYK0RmXgHsF6ivwx9SuFXEmGk
baIxMoQcha1LH71xFaWZM3E81yBPj28aQS/frwWFCTCx1xRvhf80YcMsF6N6aEfp
J5bDUMxpgjHdn2HA1eJ0LSZiNnqrPTMXr4seQS2dn26YDyuO0M4pbx7ypE+AsbWy
KXy6bJXu8Wj53ZRlPNetrfF1137LPFJEQ4RfcI3wUlYW7aloAc7SwgeQnBczFA3l
QrJJ9nVN8vr9iq1/bJ44fwdBOygLY60+Uwa/8Ls1iZXvoeYkiKQiz8xdCqPVHOIK
piLmZgJ18vGGRhBN/hdffii8Sss2xgevkpGDwPSuiJMcYB/e88krHpwZ3/QwLvwe
sH9emJv4U4dZg0ZTOeSi5W6GUmzZy8htDtfcYA7MXgnRJvdAScRzRMpZNB+a8w5N
iPcWiEiHS/lWtGmZvx6JOnI5+iOHmNdCUTMeYPSKXgN4l2qHqiyRmXb2+u2Ys4Cp
lS8wUPwMobeTK9FyeE5jgYSscsToazPaVZiL/OceoHB2J8VNg1Keo7Tl0I4e3j28
DwTJUY+1UCuzNn8hiqjra2B7HW1sTpmToTaculSxI5u1SmvP09xKlrzmwUUUwXAZ
I7vcO5Y/gpinH52ZLYdCkntAEawSGplFFa0Mh2MUNFVmQq79jui1tQZbI1qNlS91
FpjS0pwV1bqr0vnyj/OH+Uftte8z+9akEzGwlv/mOzE9GlqDKo2+RZgsD4KnKQKf
FmJfgpeUlU0TnSpPQzb5WjOfewK1rMHbdhc6hEQMmKXFoA3iqyKVsmS5hGaX2t+q
UDCzmN1UL54c+p6PxzYaB65PffyhqW8V6Ja1pV+4DVVGBUQ6ZrhdqTqJs7P/j0Ts
8lkM8zccLEr/B5ttDIZRQ0hmYG9EjkNgqSlyPkm1LYdrY9zfewAZOSYQ+HTR6bDu
schFVHROpNHonibIYeNiPSdnbSmMkKUewBdBiLHht/w25yPW0EN53Y4xuCpPXG4q
x1YCam9m0Aur861b+cwhkTzFoE44vIV40A67Un6jiuSaSWqRwOp5Jlr3YVKxHBp1
A4Gyby1a83cp7O73Osm09ey7yA7kCG2MAAgNhOFtD6J6LJ3XWiynm2hTtK4ARN7I
gw6TIjLTkoX00tHJ2vuK0dJ4gUeX3OsFKyKPPUWJXW6AVoc41x1sXmM3osBp699O
HWpiZR6UX51utllld80jdLhkqyooGfhA+IVANPKfjZyDmaOLcB0UudSbPh/ruq2d
yFhm7oVG3+2i85S+UixlC++Vaovm1lTTFkcboHpA48m3wWBQmF6CYS6eXui5Gh72
+ch/eGo5TvRw0gSQSMk8/ch43NOZSYN3ExzwNNVRqUhpJ812CrBwUjleAh5IEVuU
EcDyNj8RTSC+astxcKDd5puAKxr4XU5GX9Zll0SekGTKKcWeqySJn+ZGkWorIGvS
+XdmOMMXHkOXKUw6SfFgRi3nfXqBRl617xWeOhEgnIbBV3j0qv26AEK06VMQ1MZC
y6cwF/E5moZxyR7477K8VwUHD+0WN5oyTjxbSrNf12jGKyv89tcU2a6MPSvsYZeX
+B5uon5KZsKrXs45k2Kwu3w0Bjkeo0zM2wmj/HF5oPUTh/TJYJuEB7uWEC3ZG6r0
HYsv8ceag/yrHSZu35jIqtrDocgM3JAlFfelTc2zkgmLBHH69AfAbSQBSPdXO8/Z
40wPQu7on6AOlHY0fTw7T+hOXvtciOkkqTsyksGIsxpcwP4yDfkNUr2i562qxXH6
7f4q+VbkjlJLa3XE8KV22Inm5Jo7L8LgtSE12F4EochsuBtrIl4QYSkObUgDMF8b
IL+/mduECBccD+KvI4tY2KdaL1wRJOh0WNo60YAtzJBDca4AX4YR1CVUmTDUgpS0
TMKpudMJLi0tN9vsaJANpexFpuwWmv0/YfEHq0xx/RMfNQ92mllRhNNaeD8g46+9
PfxhUBN3gtA94xuijbiaYRv2zM0LA9V0PEZ+I2G8KmUKhvZeX7ns75PM4I0rpTPz
nIVlN/vsmfMuFafhHihCvZ6C9fDdd9RJLWAzfrfHclnWzzaCbYgOWdO/7RrDxr/k
nepL0z8m5LmFUo28bH7iYoavz7KIduLpLPSlMrlAsuwkoG+uFGHHD8oEHcmM/6YI
nypjPQ1PlhXxnYhYcaSako4zKxQRA4HixLTRQ1PdthOAgUsxrniJnIwYCPsB7ujc
kNBqK/2P67ajoFG4hua1AAaPrPMWfZTRqkAbcuA4KCMRYMZiqiKz4Z4KCPk8ycKO
RbsQCO5+FslGHfEUz6qK64I0S3i0SVz3+DxX5MJciPWFxmTcgQhLehS1sunfgTG0
Bx7WP6d9cApLqZLftYBYfdlB7ZQY/EOf7hHVFFLKOhJL0RwXuNjJy7RNSwTH4zju
DKBBPUnieCSa+Rru0ZOzK0jlZ7QA9Q2LyYwO9bzg062qj6JKRO+B9KeQU2D8ZMUx
OuAsI5V3fwmJJQeITIiDPRjZwGiBur7aKrg3gymbNtKEGkDQr/SWZ7oX4uVWHIhI
wsQ26i78BqyNmGJebF0asSS9PhZ32zL/YxUc1+Sqk9Y048OGozIaQlIsWeJ9AChI
Ino/eDwauMhu73BUF47EKQBlD5Pea+BXAay4IOxsy13RRFitQ2OJfX3kJnEP4wmb
5XqnzkCqJOURmwqWAZz21QxG9C7KbA4V4AZ10r6+pecYmZwumW2lZYoUU4MGzEYT
AE5Vl7bWZwdLEzPfAzTJmJ2/hF9E9lUZQUCk2FXHAubYJgeQtxnAtsBmCfndUz2S
rh0Rn8+pnIlkXSXFW0e0Iyn+4OShYxBghjok1bisr0U6OnX7HwnlWiupSLGFPp9l
F0rIAEdEQTyrBhyGSTVEWGWBA7GmX2RKR9v08aNhoaNOUt/ZgH4ZgYL/9wy5Iz+L
a2NCbY8XmFFO3cDGICF9nHffi05HjpZvkUVggvkviOqRw4PZCC4YVtzzOZhtaIVp
fXryWlfv5IsTiFyAW5GAvQH390mW0DJDWBq78DUlChiiF+tjLlZwbaWGdSyeK+wn
MXcg8VkuwDHq8BLA+OeBTVbZgNnoO/OBAPxQAGXagV+u4MbJd1gJuqjIgs7qQgOS
fEAJpmkdhcs4vnrE59/oaa02W+BKxQU8fGqmJ8uweYjcnD512QMhEVkdTpzDgxqo
RQD+AAkhpDyZvDhrEXrmp28/h4XIA5ISjqLECGOXBzfT/ldIHUA+ROsQdHdNkXEx
FPgwpaUCN+gokAt2r5eSWaPXNlyP8nTQx5/mXk9juujhbHRDKvQJ3DIWNBRdVKhQ
A4tCFTJwR89vvuVtJKDN0geiofdQ7n0I6taaCawtfGxjo1Cq1QPlDheEMDQRTcEm
XPNQYB9esr/Am8HcHed9xrA2eWrDtUPpDFHtW+AWKq5UFvlqgG9M/CBjN8VB0ecN
7x4QrwvJfoAPU8WvZ0QK5zctJkHRxftxmANoYkr989qCnSs3tglBTrtN3+nkvbJZ
WdxrmCADiWRVbirYKXZ8NZh471FzQT6wE1G5KzUGK4tISVrs9s1sM7CSAroZqrVh
eZMMwo5PCZ7EKt1cBGhtqwKH188sDAIOG3tyPQEdKst9uqImB+RgRF/cplP38oWA
QMs98I1VBXkG1FalzweptafYP3aCKD17OG9XsBOkE1J4m47BQhipjSxVohpLxOWR
44KgmPP78DIrGTBrmpmPMALtfdiW33kChEis3TWN+jBjyrruYkHOKCmxtqcfdvP0
nBaBAjKGBU5mtVKr1p/yw6RMTaaJWAw49W/dI8pcnpptu79AbvCZ9RPtq2M7md6P
fd3k+6v5cZNjFvM1lIsNC1tiROTL7oqUM0D4Nn02CWwZggjNGrQElcXxWj4KsvGP
utYGoUk4w5MFhgZPf8Em6PJF8VvB+NwVhzxnHfOTvQv739ocrUWZcCou/NNKDmcU
1kj0eCbVQJ4bdhD9O8pPlm1EEwDHNOMjBsM6aI/k/n+Ah+3CGQdpToV2Do/nLpyZ
ruPJ3qf0Ue9phUwjtyQqkAS5B7nIqk5mNJzsypXk+Vw5hL8dnFxxAuppSPuxa6Sq
msqK9mMhAmG4JO63B4Khs7DUFCHneMARRjnqyFrp+ekNdgr/Yx+RSObLy4wBOnH1
SXNlLWv5qJ3SLFu8gld4sFt/s0/qvi8LqJEhp9d5hThha2F90k35DFOQKhQ9bizp
7eVslbruLCzXBPKIAhmsfBTjzSOh107/7R445eYwV6PX+ToNgFIzBzi4Czj9QDJc
QEWqptZOTDXOkJ5aAbG8W9185+Dk7ug18k2rJI8MBz8MFz4PAXHh2qe3tYOyHWUH
S8SD8YwhS+ryRJB2kl4reFey2gHsQdO9VRkyKu+lPl3JByr32KVIIbloXoYF7mr5
cU/J4uZa7skcemJ0dzK0t94XQlV0DyNicwUk8O3ztD3IsrFZNmFjRuHh/9UUFil0
FW2Tdcim3COlbvV1+xL4ylkdvoHGLz4Ul5STPRSdFOa6Y0Tq6CqBcQJ6Xz96JhB2
l1kKo2vbJZTFD0+L60WrPmtlio08Ws+Tm8pgHeIXI/dwQUzXYpO88NInUw0/nxSe
+FifyL4KEgge+cZiTk8B0mbv9O8DO+ANM+lV9/mC8+oaSc/ZeBgrpc5BMiEOT0J6
DT6MgHuqGLqP0jO5CBA3qeC4JcdrxZ02vb5VvGaH1xit8p2IgBbfsRSU1WJv0YrJ
ki2vtAQGKvC8iDUGCUsYyCdpbB6G981NHYkTRKYD+t1oglsStxqxME2aIWneCWx9
m+P/4UKntsLhnnOxxKXu1+os51yY6cNPDbs8aFztPMjvOwsu3IbFYCxbyD7nFKtb
wztNoxOPOh7pJPNpTVix18oywDoofOyh+7s5g5g3OaoW58fGdBEWCoZX7ov+Mhxi
3L7R+8QzsiG+65lYRaM+WJC314x9hNdf/FtUYZtcHcEfvhLfrm1EZMyLoo+l1He8
OkEaHO4nWzMNXw3gXs8A2eroWrkswMp47rD4s7Nxi2Kfmf5fDuzCpYtC/omoC9rd
JXA/U4rFzRTwihD+qYxSWpFKXfgqQ3s0NCelqpdSMwtQyz7DWOXyBzlqG7dJcYXh
wDZewASzDH8sIfe4ZqC0b2F0skg7244s+Po3uvP2HP0JHTEP2xKMo/irocm092Ou
Dh0qAa1kNAn3KLFkt3nRdLlqB8lY9nnIIyCLqk0XRuHbh/zlNP9SEqMXEDOBdBWs
jNur19eze54JmClinjap1gX1Dy82EJuR3XdluTTBGkyCGmZfzQjA6LmC+AJczi4a
J7S8P8cKIvDqRFzPhwSZPlwCygtc/zhlixYvvGfXH4xFMKl4eGmdVkI+Oa8HR8qG
5dWobI8L5n+mp82+7FnZuWKXUadKJb8lURxuXBvZZUmxf82LncSGgpUw7zw9WI0z
rJs1E8EJ9MSx1fouWC33+M96dx9v+4WaEhRBEg0zhJU9e+vzuhRFHTvNvXQy7urd
DQ5plCtc7tekopODUCCAIOhiuvVYYYt51XEvKDyee4O2YKJhEg3jpPaEtfsHjigg
kw7xNvGEE07uchc3hcbryYp1QvAaL5hp/g3XUAIdpE8mzRx/AzDLMBVGlqTnFELJ
YyQzFJbWWtdLDT6cjq+hJCN4QXeFIRfCVdkdhDfyGR2jPlLlpeZc/u1Z8n8aC+49
9ds+zzohqLAo8w5V5CKIWBd229vVVKiKWkw6I53xf5tdru8ZLnrGbaYh3hQ/PUD4
nv6q/nj7xVQtfrRrquvaq+bWZj3ArUt2lUVJ+PBTn3yCPJotGVL2W1UGCNhC3sJ1
89PC7S5RflwZDD+dpJeOGCJRjXJ6qqN6VgI06Wg9zBAGe+kcXgVMMtl4qzHghjPX
YUyPNX0lROE4sZp572Whc3RJpXEF4ljGAgcngZN8XTMUdPNkAYBI9FVMuPscwhTq
KbAMWvwFMszSMeQe39GlQCbLP2ReGnFRsUa1weOM2VNYuUujWw+9FV4ws5LIdTQ7
jG632U5Tg7hdIWn46Sg0vm0RzFOxa881+kSf5Fr/32lu+Gcvf7f+QCbJK+Z8w7Ae
FOq8d1JpVua76AMiU8pZZPoJcGUOLoUnd6BzgS1vzUscodmkK3tw70oG9v4CwbSX
aijheFMnEtA3rhT5m77FqqP1ZREmAlkiqr+t2l/qTPFJteXj8Sl6guhlgmI3nwvV
woGD5DJKpfhG7Wo6FGziwtZFCG6um8aOAU1wdR3d7QegPKojFAJzraAkn0iTTM4t
5t6SuMguXXlg3ZPnEzdKKp896ayL5o3+4+xNwE4ZmV4YdU1SGFGXUZkNQAqcwXlF
aMJ1CWJAS5TEiNPvUKTexO8Oxdnx9A89JXH61uI/QuwSM/7yt6UqP5DnFXvk0mHJ
qrSj35A4x0Cgd7X1BKEnHGTWUHhAkFyOpe9oj3rAwKc2yjacSPFu4mIMvKI7RUYe
4Oa5fqUFRdAUMj3pH3ziLBDuSgYO0CqIhLnkKAXCzNUaFuNZFMr8JwimZ3v9Q7WZ
wqJsb1zpMcq2Scu7gOrTtL1HcrrhL4uvwqQ+zEB4KR/YFzrudxajKDNdevR5QbBC
/wTaugOvVsy64luI+pWIk8evK8w1CO80owVPftMuH1LCRC+55D/ihI3KrLYV/lzq
6j8MbuANxXKYEHLX1FmlywCipKETNdcYqoRVFGJklHO4KqXCnoS2K4m1hxkfCcQO
z0kehPBhAH9ygUcozc6/pnK5CT1Fd47Bmp4AHmswkVZ288kTiofCw169hG2FC95X
XfpNnxBBpNtwWajZEhWMhGKIM3pW0n+PwIAJUzeSFZD3uJfp7bkPjgIlZa4BiFFy
Es6chSvdRAGzqCbMTiJ7ErQPNv+qQD3faTf18kbSJTJWJEnOOzpOn7dVZy1N9F44
EgkT2rIcom5rnbD9huQMW11ui9HPhbG4XnYGuKJYAnfK7veHPJyVsacrckv4Uozm
4vX3Imt0ToflR/vSOo9GQofwbSVZtCsLSvwue/NzD3vP5UxADe+ZBY4BciFOeRLw
FkAzQmVcwYpEXswdYhoEeCsMGf5OcdJiRJ+QpgkgaSHOVRN0vdpdSMkRgPFQ5SIT
qkdF9rZiQANhLNY/DrTRYLDx96ktnMC6HUeivZ0FWOCN2LF2FvVQIsUnlMsQ4HFR
aS+bxVasAoNHyv1Rq+R0n7GBiZ2rxTHTbSAx2WaZriF8Y/FcxYFJ/l29wLbT91bm
FyeykikfM1WOJpDykxkmovy0jGJIbdfs8qAhyeaKtCCV18J2VX+5L4QX51ByrnTB
RN6X63Kz0jLRvdKDY8i0FlOYl8BylkoFxuimUsaxyfGVMr3NoyVTsF+eKzp3aWfx
Zvp0lqAgkkOiiypx/1TouUM5z3HcCAxfcXiP5mv/xux69MZ37YBMyuuhZyYeZ6zA
MTmPQmOlK2LEixZEtGdJvUCVjNgZX/TxGZ710NfdZffeyFFHt3El4G+qPnTOxIjp
x8Uuj0A9JNTLmGDKqDqz6ogStsgg0mkzm3KR0XKlOKBUqVGC+qfNF+29ltmWl0V1
o4lUb2k98MA/zJy8YdklM24kplsPG9PdGEorwyAqVJfXfS42d9FHJ8cmKSkJSI50
joFfQ4Fa9FTyLonKe72yQjTe+PIKgrvicOUsLUBv6u+XmyIrH2ub7bVLORuDBt/u
ZyRwTVH+Nmr/8w7Nl22Ej/LoFsTl9DH+q5PSu1Okg01RQAXOTGkodZpwlhmVjBel
78HluIW3pfrRsEBAyRolUC3Zy0Qfkh545hjwOo1xNEFm+79pLOCKFRIjltuJtgxW
XedV0S8UUSofUFS8Mu+COsUT468L59EfG+cqXyE000150r6WI6Jfy6bQRYrRs8ME
CitW5CgtFHKcnaxsok4hlONGYIv9gRthl1buBQVodlbhQ6C9Iau/u441ozp17i/E
z41iyv44aVxNZ/fZ8O7gCIR0Im3By5ZOPxUHfKrLfs+XGZMAWDOxqdlhhTGzMp2V
JQSKBiO1zeKz6xw19bfx+O7u4IZIEnjWw3MZoK6adcj6KN+s90R+cf7IFxP4rUhq
RaeVogpTFc+zGN5gwBqSIdywt/OzfKOCVB4PWoniclqN3AE+7dEiOdgN4FmfymcY
xPo/xkahaBKRQez29tdmKGOBzxWBW5Nfs2dje6wRDnmWCyeuZhKubGq7xOZVcndF
i0ejNVsV56ozMLAtbX3fYoQa2LTseWAFFg8lqeeHOCiP/YbymEmJVyTfIbqCRf0C
p2xEpBsj2JtaP7aKxwAi1vFEZuME00924StIrnnCnIA/lSTXI+s+JzK1i9q6375M
QTqQ5Z1+qLcIo8JyYa5vzKbQydPzairOGP7VnG7wEjFtns9IBqT98uwso6akKdSI
bG/b5O03XnMMs1a/Q+dR9RpwFKGJI0FCotmT2O7ac6mabIGIjZYbTh11ZcgrsQmm
r1R99Tf1/GNH3P417bxYnIlnY1Qr739TIJgHVswRizKuQnjBG1IjmZGGQomhBbLn
9UbHNe0HO2TtVeEvaJ1VDHXw7weUDL2sLSE5nMuz8oVFNO7ZmXp/H7HOMdZZlhOd
E+T8h2X+HqUVINbiHkUXRzBd8wx7EFrB9OpbcGq14O1pfX2JHADAPzUFFCQXHRQB
4YB7xnn24cExsU9I8GE8EEpqd2OFi/OlCkjpYhjI13C+eIf2E5LkN9cFHkEjEGJq
BCNGnroZ9CtLIzyFRA1P1+MpXJ5/U81ViAQQll2fGlfrFfeoCjG3mGc/s01gmGa9
GprwZpnaa9PDX/Zcio67/LgPm9qYMq62NZOE0YjYDv0Ml4umRIcx+mdAjJI71GJ6
KtBx87DGj1QGoek9zOrC3DzQANwKaUQjkJ5qd4lukgS6MwyI5e4VmwWwsNUb7hud
rjyUmKXod5gjWpkzef+h6xWGWRcpemIU/+gH6NtObhjMCVgg0onA1iAHpP69e/d0
CBbC/NOVRJLMD80PhHisq6sf3DNIRVo7GGIBz6QN/cjFAj973dUyc2SuZLqHNxrL
lz4J6nvvTmRH+TWFdG0FjzUuezQ588ny6EHbAE5+Q9j6yTn+96RZob0OnbodLrVB
WtD3RG66rEKh65QOLhkQdlAA83SvbuWsm1sGXc70naO3tDCa+oMdNaHxYKt0ER/T
EAWx38a5cWLO0r7qd2VlOrJbOjyyoSqHt8YsQd3rdn+JrHiQMayCjnLiwRieKAXj
B9N/SyIbmFcktt7GlG5+kZ1pZLTkJ8pES5dHKFO/IQTC9qCHZKDvY+onW3bOa05x
4bvcDScpTc4VGB8xrM02DQOL4m++AKSytULxVmqbqouvE5yFcRnfbZrFiorPb5Fo
YXY5innjuAc/7RTR9hd6q+f4NBmZb3vN9ZT+JEtfRISf009wokJAGD6zKxkIFw9X
JZhUS6LAjSasKrb6B8iN/Lk+RSS5fxjk/q1fHsc4Ce6TqCMRo8/Zopa2OWNBSmtF
3DvuDeK2DHszJvpzjvIZpJdXAUc9IysGcNLFJfvMP8nlc39sPMLlzwEzYCO9Lbgx
hP7DRhNCE8+s0WQngUKpYO4gMhkWjyXxTZkeldG5sIKDP/VcG50RnfPxcTEfvLHC
xFtajWpGoXH8GrMrAxSQRi5V7X/NykfRDk5zY20GEiW4xEPjvrqeA84wE9kI0tV4
zrxZ46dawwTdsoOsk/r02MpYFyE7ZhHJyn+flr/aLLrPhxrWiufyhaSZ1Du7ApQB
wXPbPBrc8SOchazK/bZ7iz1J1b+KaHNvxpevFJz36s6L335uCB56hEbWs/72D7RR
SPYgvwmbCv50dEKB7DqI1KgmR8w7HzzhwrCvesCyZ6gHeiHQc7w4bgSy494ILvln
0LZeoYv/f67DrugGs4gIv9NWOiaqOW/UCiDh6S7MNmLWwhUqbPZ8X+Uy9mJTl+7S
6wtNqNEOCeCoBpE5TBCeSFmBCVKilXsKPoxS2M0B5ABTnfrTQCl1SyJbFjyAco4O
0qGdZHJc+8GwFjwfG5xWur/uujPUQnzPxUNqwQtjLTvXTWW4y6Ulw7S8p6goUgif
FhYqZk/Kp/UdngQoVhCBby5BPHNLX9BIs9Pjlk9SKdHxoM20jVA9zVVyM2Mw+H8q
euIoTQub05i6MOW+PXIoeQQD9O98yCCp2iHXJ6umir2uKxkKbVMEBpJzQJHLOXtN
by8qTXxIrihPiUHGKKOaOH2cdlmtwO1jTJU8pRDM0Lqejf6ixkvVsgpUJOaxXlD5
x14+NczRVyMwNhnc1kHxgqAUaQe85egRPVDP+ABtQXIqau5oIouejHRcGUTI1fLY
vzK4jfX2lT3aVZx4vQEm5mctXUeLXPQY5GW4LUMKR43AyeQXbsYseR6RD2+6MIxk
bRS3bnwPkyTQA76oDSd31zUtrE6RmeRMXUZ2c5c75NXnvAqxMtK/jNUAzoIzlErw
4GLnk0jNZqF4UbHHW8hZcUWwrNlS8PuDybIY61sHqBxePdAEEhQUHlaa6dRw+Cw5
rNy1Oppc/gLmvgebhLcuqzXW7bHzbEBV2FP/8t97TYNdaeRHMK4tKJ7WPhRCaP3V
f8zLRNCFEATkRPP4YufDmd7/DoT9P93GXknZcXdgBch1fddyGBTfov3OtWlZK6ts
A389PGKWv9agWHFIVsf1yoi/vPQ5I77tzsCE8oZ/SG88mZxC4D9hpwJwwToVUP7P
4Pq5K7pxEeaEI0unG2a3u6LMySMPFLDAGxR3qM/HetvyDQMB88fnSefIFt0MJMp3
Ab7ZLXRAGmuM09kob3PM1haL9BEs4DKhw6Ez6RQWnako+mfF+u1tqjY+H0H4bR4i
ZP461G9prCqEsga6nLPKaY52pDB0c3r+hcYuMrVT6VcYAohm6bgNcgEj01sarMWt
VWKEQCuwPyXUBJLEui22soHzkCYjj3afGx0KxECSIjYqA6TGSOat24SqV9uDwmQF
4RgnOtrQaYHLhCrypaqOg56jGhsf9pd1l/KghMTzTKfeSa2PHxGWsnpM0uGpJKsj
LScq3rnv+Mf4QLXpy7ACI7Y1QLaLmkHIF/VBaEoYC/JjzC7ivMDoPwsxAndyNY6Y
wNyPQFu22BWY+AyBk8moQex0mPSRR8xpdidnWUdA4g6SaxjoWvmKWihVrpGfHuAP
d2EFH5MVtH7lKA9PlbuD8wa6VeAv+Hn02ooPGuLVJh6tfuGCirWP1/GboqYni3Lr
T1ily4rWivxl/jxsbiyaTsywBYPj+wADRLJpZCN9B6Y6nGyW6DjHCrIgR/TzheQd
OUOWrNrRg0zc6WrWUGh4MQsPCIN4qKxeenf5zrHwekhmxja7hewm/ctQRD7fvAya
YT9akF/aF2gjBszf/Q5BV553CtxL3utLmPxbwBrzMNpqgZxj3wj+UytBC6YG5APD
luJIiaCtnoZXLBO7jgZqutZF5xULEgEwd5m+xMgJMmi609AVau3tpoQp2IQ1/xS3
Xwjz4s8uc0KooBeA4lh4qPcYVCMr58nWCx3xVjvIFexzUM8xQ1njf8iD3KZru8V2
RseRHFQovZaStEStXbCrMv68PwrmFDgubV28C1+QWgJ8YfC1G/77d87Ne2ShZto3
KttdpUepRtF1qXqMGgcHjadol6FhM9IEWjZ165ykhJ4EdYDMVMPRPlf6RZDtw6LF
/PW5y3wbLGKqhPHeCvScfpzjKsdXJj1sLfGseqo0OrjFB6bxTWewARe7kR+4/xZq
fMbL+vkWIhprSpcvDfThvGW/WGSN6Jm6+lv0XIG/H8T9Bqnq6K55eeXrFJllfLB4
70nkMavsRoI6LTq91VOYBzLRCcb3IYqa3Eq/ivMO7LgVG/Ijf83FYJuey3ualTGg
0Yix6RNV7MuvQmOlfIiQ0EyPX3YRtu86WrnCxm1Gasfo6tHuSmCWL7zn3tkrJ+1f
Li5YH/+QKRZN84XuAMM8pFBPy+Eu+ZXQX4U0Tc6Xjo2nZk1S+a5cfoOiVo0Z5fIN
4i9mb3Bdrc3ak1CjbqB5joZ/vxyjUmcMYjHzEqwTyoE0ppr3IqBtPO4Ngt2FjN74
7VdXse359LstUA6WqS1XPGuJPTqZg10acAjxRuZaW64T6kjg01/E/iiGWUi8Z65Q
ug5JvkEJpJ1zafVuUuP0ljsCLjsAWgSGMLWoG0Z1R5iQexTCYBcLDnyCIsYyiS4N
teHUiNOQtrTvphmU3f/sYM1r3XGfoNaktiE/TaZrUJBawAF0qX9KMjDCuqn0IYUa
os49Mv9EL4l44fHb6ZeQUV+j+lp0vcKKmky3IqDCCcmTY039xrDOO6/UzKt+HRbk
SFYDa3JlKjaBr8cEb00EhBh3DC8otGofM+7qokVS0WkhlDqe3fs2P+cS6nx6ilLG
yBlqHvle3BwPdbcnFSRz/k17turG8kGSqjJLVr57ALjumR2babe2RX+w2wKEkbAL
rKvlzPbuyocrHpDCXy9/HCvDMJtCOvBjFyd1ddaAUcaphDAdj10OtpDZ1tuxpKjy
/E5xK34KtU631Yv287XpQ/BqZeMq9qWLEuuAWGHz7vXL04c83ykZLlE5ND5zqK0W
JAQDSw+F/xualFJKAPNoDJ9WeP5gDO0FuSeB9as9vsRyN6/aNc+ZQQ43gI6NGyGo
wdRIgospItrqwbajmT0kmrP5RqjMHoJ/PDTWHQCcBDGIAec1sRKfwt0zGnV1zU/0
zl1p/ku4KwouryBqgfpC4N/fLLMWs+nl0ZJujwrKrbvW/kbo5hRuSwdNSkBbmyAv
TBcJfMY3A17/2KYOfHTyi1fZ/pvQpHTCtDXOQaCiW/WVCMYKWjb3y5cqweDV0S/T
VfWMlqVMyTZ6J2G8JINAhIZ01e30kXgGgngdxjvcE0XXINxx8Xb+69DThVTvqW7i
mwoeLNvd0UJmKUSV7kb74XB3cH+qUgQVLXQq41AuUtPew21kgFXcSDaeVZklkgTK
eSB6VDpoQxZy06wSr+tvqhEfmb1+veenPWjVbvComgNhukVZU+xDwDToBRXc/i76
rRAJDgo0P1pVz6MIlSMdyW4WQQjMJoGpuonDWNGerLMTwA6CfAV5VqEZIqXakJea
wwZul0uCFVAiYvlLMji6P17wA1pPu/yxihUDdxAOO0lL3NxTimcicFQvqeBEMsRx
VlsNyF/RxiecKIRG6If53dUSfiHfVxSfh+VN5m/WaR9u9RPulJdxqHg0KSVeV3Fk
bs3OuSCA2udyM6XVUueo7DYLUFFZ0oISz/ELv1mbTkezSAsN/44BirjyZdb4lprh
mLAWvXIEImwn+TTKznur5zuJPbvSC/03NmThs3ontB4=
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
EqX0lGpCzwnaVRh+Wi8LxSWBLwaPltRTpfZOz6g4xYPEt4ApTE8dy8ULQPT1DSJX
78aaXtIKVRY5pYIV2kO5tKvZ6XV+hxodbwnMffq8tNoo5fhvSZVDnZlsHZic3jor
mvmY1MeEk1FqqvFVCcwKRr/i+Kv4g1ObHXx16W4R+T1y9mS1bymYiAJESWYDCeOx
tryH/tqQR1g6+bLBUHBIu+nBLNsSQmKxlnTlSDKCtzE/5A0f45v7aS6ZN60TdYQ5
CJ1Lb1ChLmBJfD2O4DTgDnVjfvB1/1Lrr7kq+CqFAmwabP6AFE3e6OdEMX1LSwUl
UtfePX9mNvX1ahqvHe0pJQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 656 )
`pragma protect data_block
ojsMysXl34+aVGQllEUQ4xEAFdk2i78Nzn1dojEq+f5Z04Otz6pwlUgSXrothNzN
j0CvMnIV6d3ElZimaUhGDWPOvbiypM9hh6zaGPiXXfOJuqL80fnRnxA8KEkDJuY4
fqSwiLOkQ415onWm8F03nzHGkqlprHhlngGjlg3TFwHqqFscXDutXksjkjDtsUF0
s+aCx91u2AYZbe7+I2HYBuiiJH66ehE3v3DyefiTuNnBdHF04mQTIWPafNIOYfpX
cenK7ia73V42wfWV262+VExaeI0z5E+Mycxf1aaXkGUojdHdtZF4tj3OrYFcE6dO
/PiJY7qZqUr9I+aEycuMlrubQf1hmptPsAzSH3/iJheKUv6nrNzugM1lThEvGxK4
A+p7dbojyYEM8wM3HvLeetUauIup8s/LwJ8obNN7VllX2rvmIfj0+dy6n1Rvqd0O
SVv89AWtIzhBAgKdQlqz6TEvNx/DdYAg3e7hZ5i0RHGGrR/znWZa/WteAxEQuyDh
K2ctQEITOWfzbH79M2h+VDSM3m4V+KtouCZ3th+v8GVIRN1PpzAn+N2HzdbEm5Cf
8eJCwSZaFh6bCtu4yGFoPBnwx9ULklKJzjvNyoU7UjLVe6nGGGIaEY1RNJQDObYp
RQ3G5tE/GEywtrz7CX0DtrpAWY6PNiGZ0rRtJFbBnWxJ6/Ae+v/Pbc9CcANPnCIW
6yWqPdrZVqdHliaST7SF1QlgqjL23SjsGczrlpaehp07QNU81E5Dofm/WIRkKc06
RQNZReBW7yQInYZ/H07Q1YVdnJokyaosIKcc/Tx3uOzM8AXvs9PwgKuFY/FnP7tH
HZaz8P/9cJnqNhRHdaNDpf66ejoueBS28AkZr+kIOR0=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
I88BHzUbomNe+fof2+tf3Aoq/5QVmOBt0r0uGHByK5WP+FlogxmHFKCY0/6CMrX1
Jc4wekjA6ET90Fqn79yCiqorPIvuLUDi/S/hsJMN2WUEHu1Z6nXoRBsbjaXSIYPX
X1FxbvHxjB2//p0SMgiLdFLk3lt2mhiJlph0h9Q7ulpzZHFL9WxkM7Ng8GJLy5XL
QcapIV1q1do7jKGNNa0TpW7RZeLTlMqgJE8cBMLQtNVOlHFnOW7MNDSWDBj12EbM
2en6/WkRmlrRSxyOivc/V1LUfMHeG4DobmJAM0p6vNg6ui476HHGmqNBJVOB7vt5
ZwttGRglRGEAUMMmL5I/Fw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 13024 )
`pragma protect data_block
LnSRUBxRvBCKXKrg65s8YljQvJDtXuRolm7NEeRSPmhVniYkFugZaVZnSHAk4Ov+
gRYlH50JtJC73Nqg+W3Z2CVyjxG1YC1rhQMR8WuJTbu/Hj5r4597l2tm+xy627eN
7RJkwdaETe7pR/OFzFWNI48qkfqzL34zdE7JZNiBI2L8fZKcj4O0kaZqgDmJ8EeY
FOJYn4fFhi5EUpbkGVt8dE/w8/TACwpB76xkftb0L6neT5Enc2j245OPHLHmproI
sQScH97+MSDhKEtozTXBBoPDcwv0/M9h1iwvHq7DxxQrCMaRbxKZ3HelOFzJf65G
PCo5MeUJ2vrlpl1iOo6EOGgtwAuK0ygpaEctG2ee1+k59Fo76VpUXzLZn4i9Eo7P
YlrXjAFcE+ohknb14VY0ev0qkryTjb2bfu1Ua5mwB7MNNM2FalmH+2LPDlMJkY7F
P68Cf7S24pRpleRvkxnce8TxQYUNLD5XV/jwVbdgtBNGgj4WnBBaTXyOJaCul+Zj
F9Lrn/Oa3HlGqmAy8WzCcbOYx0gjd63q0+zEMQcLthRtwYEpRFT8qHhE1egBujXl
A/ZGvrZWwmY0hcmRW1PneErk6sXq53FkselGCUYFP/tXNKBbMTmILpAYVqdqltZY
/WZrx/VNJQRgJYh5RXeMHaqEMuHIJ2S7Z+z6p3p/jQg7miRPUk0LkKVRsx/of+4b
E78Ea7kxCgd429HQoYz0C3jo3PH1kbApNA8tYPKfoJbvpFvQiMKofZyS6p1vhLJq
iZEGt6bNnMOFL5dxGs4Ho6O6bQlzRbYm+1cXiNzQAQ8YKvKmivfrYdjqVh0RKPbV
sCSJgzYsoKYfOtyZk/GrHXS7JX3tXsrWpqx+q5tvhrkbEQsfjQrdFDOHCBtEdR0F
IXJ13bw3ik1nX9BKR6aMq1oR52CF3Mcsnzj4lt3gCeqeV7phn0k8ntvIrLm2YTXp
oWHUjAmT1X2wNEugpLuOu6Oh9LqBA4TQUgd7R0SKaeXr0OsrF+Q8LVdz7r2gHtz6
bjnXkVx3iA1yAUYb9emt8SezSUZcioGJKlK40SoD5n0xEQHMU0jJhKet6fu555Hz
tFIpLwejq3meitx7+pRhcyLU6CstZ1Laq14PQ8kR7I9kzUUimBw6AJoZrytO5cGq
gP/UbHWbL3gg2CGKLQTIymtmA8jWHfQ2d9UKymIXUW2lmXmF43Vgo5Pg+wCW/aSJ
xzVyHLVAidE3V4zh9KLHmlCb7fLdtpySYiTQEjsVaKBteD51ijp1V+ZfGAsL6OgJ
VCPblpKbBxmIDSfqtc43BGZUeyF1RnZFXBErgTzI7kVKRK+DnkDcj2qiPsKFia4i
QKY1fD+PbUhA4P2jmJx15uCal336hf2dF7qYPLOjp3/uzwRwDOCzAdqM/8QcE3Bx
OYe/l37NmrQe1EDj/rZbwjFN4HwM1nobdBn9eCcAW+VbXVMSnwmcYaQy7iEwSP8N
DOVSxgsTcSXffflaKkR+ujF/8L5rfm7v1l6LH/CyENtD8KBBQLPB+YnOrgsLbPIU
S7cL7klenhUFtHoCT/MWRV8bZzMDdKf7gey/0saxo/xKIziABoMUWa3CKa9U8aak
Cr78LNxLwHecfLbrm6rXn0UnvquGCJ55zwZsWaZGL4IN2h7hR+oBlhVgnkl9XOj/
+N9xlZCkK2Yl8rT11s7pLE3fWgi27vsm5TCgjlWmG7wiqyQ/MkIy2KiFs3GKFWyy
yrcma8ZqAfePglfNy1m++L0eab9JINvWkoKHntWBLdJvueFjHjBs7KlsQKRiYMfk
tPaXmHPQOptq3G8QbcMjAsfySYOpJkIAaVPW3ZoMQVHNT0uUo8Qjcb8+cU639AbL
eeG0ZmT91vzjCXO2XcGqyC6V20+YAJj8KGmxmdCQz2tQ8khzxsXO8G2yBMR2FzSJ
/aiQMATHafTzR0wAvk84xFQwjxA4c9+uM0VOqevEGZR6Ri17WOP+ZmXvjgO/pTq5
/rzYtK0pO9ujLcUn44qlM2l8jJcjLeXRC62vvsoRiZ7auqZEt30h+xYZxm8Ha84O
TekkZLpMAJQCQLTqS/jJV2hW48lWDpfr3wsDg008K4B8Y7DjEQW2bPwfS+uw8CwN
DB4cMMGsITUWpPV0Qo7DNLzLdbLSQOeQR3M0CfnZtTQ9zLuzGfBi8IBY2YBwbksq
rDHYa3138qbfagXbD4qGQUzT6BQRwez7Uxlmswt7epE38CGsqtSUathj3uJCuvoo
Yaf4EiCFaTkoR/3Y3STQWVWX27ItGSI+yPK/24jBFXVd8dYTI/6jBQNrJqr/vbs0
pQIV1GtEGR11G4EtP5CPRRgbNIn6O7XMZzGm0rNbPD9agAoQmlnpWpbjia09niJi
H0w04jQzavTqAwdjor2jx1XW+8Zb8Bxsw6HBXva3LpJ6dMGBM6/l9cyDB83DcLTW
6CIzDh6T38dk9Q+v7Y1oEjbOuo/mL4CrAyOOeQO5csLNL62zSKTJvzF/2tr9Jpmu
dn5nc5QgVxDRX+1+dRdturreTxf2w1K2AFNsFsWRB1BgNshoH+3NwDcYY3kVV2lr
GzoZdkqQ6EuI7IDY3Vb2Kc5BTSjtdr2bj+T3GpOaU/13U2laKXPStCmLZ/6o74lr
/TUJ8NoycJxWgTzuTSiFeLj+81rtlX3L27FnZpYKyRASg/2Wox4l/8qGKJYTieTu
5pADzQ/qmMhe+4kttZc793dsdeES0e6BcODxpkwJy36pTEGXHQCsT4Add5TzsyYI
CukjC3/lFMyRYvVHqjpR4qFFnofJng2Ihy7a3ThIaSp3HDWbmWQqGg+GCRNrPA8c
+ugyoQrrMwb+jdkLA9RnG1pcm8jYaXqLo1WqF3cjQd1uSK7v5OB8qkDy7HviZ46O
eMWEal91qpF1o6F52rjRn+tSNKrnMgbSFVysvHqt134WT1gedaGdYxPT1MRutWR/
zsiCYyV8DTV4yBi7KQj8l0pa8uih+uElM0SK9y/39GGVKaOrCF+j+ProwqmT5BIZ
dSwdqbXi7RUNkWHiWZ4Dnf8gUQpjkRgcty0I8PmCayFWPtRlNr4I8psRWXnqNAfH
m8ZJf1GeYs1/X/kgvpP3o5myXpNeVDsw7AYOWGVJeEBuBcvuk7ZU8Y57Wji8ErZo
PhFrMay0OhHLmJFY7Qlrc6gCXecSxjxgAQB+tAJEZjQVu30jYt9LjSSBg4l9tCwm
WSl0kW7bsA6N3vQH6y+PUu0Ik+I8wZ2c6WwLNcS2NwooUAAderqRV5lPLCDtaAVX
1AoxLjmti94o6exRq6SiHjNgjy326y8B+dRAbt6ulmBgk4FzPfcAdk5hAavGuaPP
DQjTjhZo/msyYVS9G7XNqYM8g9zPyWUaMsf7yeyxy0ZNoq6NvHmhwwQwYUh1BUZ/
mVdh2pUbkbZRuUwKp6yMrVemV4nxmFYLRG7Fgqe5r3AseKRTx7esVG1bimntfVlV
5u5fvmn+RVEli9liasdxPZoBTrZ6NmdxXoiGx064ApiqyBd94fl6TytOmCVxKoXW
KVnsfIpPSuAQRuTqS4PEHiwO3bpvEwxTYqhwfxJ6VPmWgq4t4RpwwsoBjDHEZSrU
jjoh6+6sSVhmfE5tjn1AMRkCz9zCIvR3xFFVFQMdv2OJh14YgX5LMuJH94Yd2oEF
JEYa7d6E0HQAuxHUEKYzfSj+5sDZHe/bwR1iClFPO1QxREyS/nwmHFwRACv7wWQy
aUrE7ooAPlMPU5YwAR+JExXcX0SNfD57lQZf8396JfycgbgkkA44TMcrcrXRXADV
zO+I1dlX2bNrV4fKNzuNFuaSOwE9s+oej7KLhZPfh4/I4h3aA4M4TO5Hui18lDra
3d5YU52ZMukBUN05VfkwOMFodXKTh/4d0Zwx9xBFIe8Mc5xu0Q7GvO4/k/TezRPk
Ax+1lsR41Lb/Ekwf4Pdx3nyiO0VnzPi3B8p7lANH8RgccI69c6H4hBxq4eqXGGHe
1Pc/Z1PmrYqPo8eAdtnTkHP5H5Ei9u9A23WUakM+jXPFgLjvyjIOS+K0rKhw6Z6j
zOK3EBweLkqcnt6ZUxvXuYh1y6VulK+WAf8+hvNSYPzeL8aQRH8fFPr8z0jRHRJf
C1T+TiV5KIdXtas4YQ0yt/tD2pQwJJkZL02qbD3ZG7HKOEZlcA4gEVSx1rMXAOxy
txG3zZjunXO2jJgipvUkIcJA//eBJTbUB0R5WByyceCZXO9kedYPfu7pp6dgMT3a
rcLvvCKPBZDH4kcYSDM6igp+UB2Prm1DlCG6CLOPIOBu67wTjcINs5TN8b+4ssTB
2MBhcRVR3aO9eFKKYrx89L3GoksaLdWoEKgn6DWCApFSaxfq8TJzVTITEa02Qvr0
Ftiblud6LHbCc6QorxoctWoPRFAv+tFvN3+E/C+TLC6PnQWJ+jXAr1TX1PnKb9Ck
iUEpvi1tdN/cB3US6Lk7e1zZQpjwjJQV3WtfgI+tD5uIvFxy4zG0zvE+Ee3LfQEh
VdxrxFdER7PCn1vHkrDfruNOkVwJVJseewWMS+HAt3bp9Nq2POCyqp/dq+mYucG1
PtxbXWfeGNQHn/ygUx9C4UAemEAwKGH9BpHsEfVwYj1dyPKYLGxeLw3qtpDTYPnm
GXVpqMKMST+KXnOh8hxPQkc2oBU2BoOFRQKU9mB7MvPnESo7yKE7AaLkv7sst6Xg
iJRnCHMBLqW+GaoxC1f4HePfzBkswEpsOIdDlVfK8HYWpG+0RJXlyVhamug+1cTk
cHThQyMhKbYVqXuuEp4uV8cYEd9img89SYh4vKIbPbv8SOZLa/SHkvDyN3vxM+pm
5WQf6UNdcU2HH+iUZVyEeXJ5Idu7W6h9vO72UOJMYN5d8pLMClLiV6qXtINgtPdg
ymD0iM7hO01UWDBisPpUBH6RDv3cznfuwwtBX1JKn7s5TrTsPDbWirwtx1XCxriH
tjvpysp54qBNS7eRpqK/OG3L0wrBjN6Qhchw0Bx+z3fcyjaQGJs8W4ERTmC5KYJ/
2OgAg2ej3TDKJ32bNDXIRPkcKfSr6HKJHlRGe7vQRGKoHEGEWTQhT/xRY2Y3B4ZS
xTNe1lCK5OFFnaXruYrwEcCeFiBPjo/PWFAtWF7mjZkrYvjTVUSOuQWUeq8cuTvK
ZVzwGCLM8HmJbnq5UipMiPmj+EpCIccEILYm62NveBMdLpWqrmY6t1rmWvdsGlIg
Q0j2tXSRGFU2dwf9CT2/TH0nyz9a83bgA8whKgCB5P3dpCXdEfkzmHVJGbaHhBxq
/M34c0ymxUq0mbo0KuQSr4woaeSys9zQhL2VV4JqeaopjZ4KgeVamX9dFU5wy+55
EH0DgusCrnuuTHT0LHCErv7nDgEqr2LDnXIHPidhbGAV0AUEdUTV6YgPLyVm8rtl
TwDcRxQmjh14yqS8B4vN/nyKT0DBO4bdYyZdYflSfToofZTYNMAwx8Gu9YKqmlZW
SG2hZQB7+hCqMNAJMrW0Jo9CuEJa1fw9fkyI6RW9x/++j8p/phIaI2cNHazPwDQk
rbLd4DFqFk/lpiXPrGIgmQkd6NeJDsA9Ypq26+/bDwQ6wyVvkcJ+xhhKMrQCojsY
JpHkgR7qXrhQ063KCrtcyNgkZKTb7MpXER0LJVm6bE8NsrPbDlamYHKueclhwwCU
Wgfpwiaw2NqaAKgBImHr0aMvfMJNsRSVSyPNVGjKOo9Rg9QjSNnruJCPmXbHiVPc
RQhuXwvy67XfWwg5CQMI1KAOT+hd0KJ6SCHUo/eBkqQIBrYES3LGwS4CV+7T/FTc
opYNDTWOYuS8GT898a72oiP4My2YDWLdBGMgyFDzjSwiTgRywPTKOOxr137mOYJl
ptKTujBoutMxUapKWevybOPbnEOvGAgNemakrmdyYQyUDLc2boD269js6etwChhw
C+FmySd+OQT3qQWULE4sBsuZXeqJL43cmQV5ckwZxdDHJUyHr7RiFdexmxh2bHuI
odNydeoxk50z45wSsv4kdrvLEUg6erzdbwCaJULoz7FT7tNTFzmu7xEN8KHDGiNx
hGxn/mMWV6IBU8SXoGe4CUwJKBtehjJ9OTF+LQ8JZPlbSxrAwJglcHdGXXVYsdXH
jfSYJFu2nv3kpSVhC6/loxZytdw7u5bFyzsPn8EKKOrt2LgUIXxxKAJBSyO/JhRI
wp5CCVsR5gW4byPqoMQfiWHqyGkkWOjyNdhkbUyv2hcts1/GI6vTljlDabj/rymF
ID/vMgycR3+24XHhzIoLG9e4bQR4CMnb56YJ4HraI0LZweMz0jFCkI/AlIi0DFPM
BtZbqrGVdsdijX17sRBaPeCTvgF6vY6no2DiFjyg59dYA6W1AcLZ4l/AS5pjcbFW
WXpG70nWrREKi4M9aMc1XMdNNPOGvBTdYz1K2/ajbpyMDAFT0iEW3NdQsz66VJWW
8Kjaenbxi589ye3824i2o5ech/CzgKT2eT9XdQb+KokLkSxMIximIN/C6u0IM4fZ
voxVxy6DEuVK0xAKU5/72neV7FNsEnqPkhgXXq1SZJNcIv4s+NEaq7c1Erv2io/a
zc7ZhWNNG22j4T7cz7eyM+HgY+xKaeYmBekiMCBbfwu3QO2DkeHCjHbFhJXmTNl4
wSx0HXFvxidYOsLf53M3BrzSzH5CnDZnCuaHzkT1XoGpc9UwRPf4X7pb8MPW/zE2
5dtCVz7Fk7xCcfUgNFmjdbH9aMKfft//cK9K9ihQEI2X2jyNT7HWbTTaDGKhYQLA
U4j7H8cWWOm9y1ebbMUoJM+Nn+6P06B4zZepZ4JYpGaKxjDoRK7wc4xOfHv7GK0O
Z2K0rr26f6JEhpP96tHaKRcDp/uYk1Mt27S3WOmEEioVtWRSI5avy8QwBpylxhf+
FOZ7n2dBeHLpN5aTHH/YFiXZOPZb7VfTRs2sdwLJCq2YFL/kDpzdZt1zy6nVPylK
UyOEn8e+/XcOFNd4oVotvrJps7yJYE3tzNLRGpXEAwhCu4Stu5TDaVlAOcnXBdmU
aiBlsiaZSGDDPMAC3BaepHHiLQBKSicD7bTNh7agA6JCK0bIQJc/EZ3mPgW3ucDs
UTtAUUCw1SlGAkaDkAmTAuqB2XI0AiGCo7xlM3u+ZkZvW+ex0AWer1JQLGGYEtMJ
xISR1+Dwc8hbN4xmX2BmJeLlYvX8DPSAbwngs8YF0o1fvDTZZQNKQo9JB/absLnd
J6Pw8c1jxcxkkqJpuMLSRF6b7l2H859vRgDs1l7JLbZCk1/UJA43FqgskiVWS6o2
iCBYzMc1elFurw/qq1C2GktPzMZIvODmHSCwtnL5sOtLHPcGc4g4f16Cbzkz3lRS
8sCL3PMl/GUFqdJbIbAyKj5Cz/19dQXEt5yBBvOhUWWi+2lX0QF8FJetlL1HDJ0P
sNfHbgcmJ1/iJczA/tOedaI9pDegKF/ACSWsBb9FW/HCTwGxJvulbtCMwR+WapXu
z1PRGTt6pOidVosHWjZyDT5cB7tJ8I9UIrANcNbAlvT6KMhw8Bte1a0R25jiQfOJ
A/CXbbptkPFuYHipdMqfPgzT5KPB+aChoJw/PVdGfmHAxvNkgjn7Yvpc2cQBfxcE
7/OSzsBLi5iepqwwK1j0G89w89S3FrsLQT2wAC0U9s1OCbbub6oxrtVASEhskNpL
xe6m8MmZvAuR0GKqsDtyF6feCJJaoJunO/JlGQZQwXbHm26zIwVcQb+DDKNEixLn
Ea665UkLMrCeSykFEgsnabG73kkLUepI++V5z6JSxHB5KTaMkUYMEYcuGH5RxIgO
YnAaZZ3K6Vnz6YoFsZxyhONYFlSXEol5aqu94pkZGjN2coUXBTUHIBIRdVlriGOW
fhsOxFm98tWSP++j3FygcoNIrKjHcC5oPJ7UDQ090xQIzWdsWmQO6+XKqeT3KZyn
m2WFpeEUfs8gO2s+v2QqAnZesQcVGGH0rj6yfkQKQ6tZ/Hmo05moZ4+f/hxBggev
WBcRFAC3lzovAp5CF0aGSlCR4dYWFJDKx8g5eAuqsoTVodqSOdv2UeM3esk8b8Mu
qtWwbWJWwXsa9qlEW3WYnatRDskF5CuhMdrkOY64HEbR4c4q2eyGTTGh7Nt9IGFi
nH4yJhwHySFub1kkvbByMY3YO4jEWEts7uq+ergyCRJ8HsaxgbYiG02lelSemqCG
ym+VmCMuei1ycPRwe+GNlDIyYvnxQa3S8KcpkFxLkGLFCwEa8jcHG4dkq/0O0Uk6
frIdlL0wveCwpyCAz9uRCj4A1k/TexhIzhBxa2m8GeAFRzwH3npIo4QX91MWzqdD
RxaF3R9lxbMSsNTgkdKJCWnIuxJSvFtqN9iUj+Eiu41+uKd1jwqTa1JPU510k/On
j9SdjIgiwipNUZtI81KxewWWNQ0s2YLU9pH/ObO0EJGnX6jtuiwbH4IaiWyH9znp
cXLdvcC1OloTlTT62oXNObxbGa+qtgxwdeRuJVPXbYMaqEo+qurZhGrygMChJsna
qBLerHZm7lYypWCJEotDVtKnSgctJHzETsOP7JJBE2ZuCx8BDCtoZfGF17GHAnSA
6Axd7iGNFy8TcPJdYrRISEj+sHMlROc8t9Spn51s78A2NhSmZ2pS8uk4R7Y0iMKC
QTtUSb/MWpY6CgH0t0ONz4KnugHfn+BhsvnyRCrPeI90sX/U4CwYkxA8GSm+kv3A
6eeKQKzcrhGwOslvQbmiVPPQJ8CvpIuOvEvjnxNIME5i11HmGRrdobO2hdbnUKOo
dJR5FNo27bBysbxAn0j9h0qwDYJmVuAoscjmCkZzZF6Yqa08BMUL2foKJvntxKvJ
ZYnbwHLmri0GR4jcQIoiHs7KALysUyNwaxRBFwniigCnjkflK+9/bR+5oBaHGUX/
Le8BrRhONU649LpZmxOUsl0zH6CkQObHQBkihExjmJ33TTl+8yBho63mKYfFX+kl
J1c7r7j8I785bKZn41w44ubyVDBeo9OBpj5U6c4YoMZJVwOEgxpoyH395SdUMDk3
tWVZWKKlxGnUGEL69DDyRXZo+J8vuR9hJrv3JoVWAZva/X0kQZZoPvV3DIa02wDi
mISIwmA38JFSwzs0VJTscFpKoMYMSi6L5dfX97lqFmjYw9wgYD6h7gE62zkw0ZQB
tWCYLOFNJQhmlCdUm5w8xAAJ0/csKbSMgsREYPwM8OHKvgqEOEGYvpOOhVKTRA2e
q9qDG4dUO1gRerTdDncFgDQ+IgBkUboJPlorxFrMzbq9DIZUj0BY5+tvlbwT6pBJ
vWbxixJDKhvBa6Bnu33o8jUR0QDlBEuJNQ42v8BYaaGjRsqK2LaNgeujgTgSIJHM
mFP2nO5Zmzypm0AL6izZbqwu9bdEFgDmXup0xOUZq2guaBx11TNC9+S3KydLudJj
Oji4uqE4EwOsU9d9qJt9Wu0lLAHXDdhGXUGZj47uEiQtT8g7WXZCCSmpvR/fvDk+
0XO1YYB/UnRyvgkB/05XLulASgh5K4H0iaM3emHRoiYaZeQjR2fSVoqONWa2VwRD
9z420FNEHH9LpiaKsl1vBggA0A8fW5m3awsYiFYZHmy0BZIQ0kMi3UHliRKPQeKH
4H8XtHoi7qL68dl+dC/Xhcm/IDoVtuUe2Sx5tukrDGaXNdzyJBqgFZzLwqg3zcuy
E647uek0hudqpq1i3vbA/Jtcq2A7FtMRmo8eKss+RqZun0L1xKi55dLQykxkD987
xs6EQdZ/6MJMl5K6/WbGNT36iffmpsSx/0esSrTqAKk5DoHedZp+AqV6SFVjQkHn
m6LgBk5t+2iS9Ywm+3yNwhPANbXe2P15fSIqCCia6EVTbrtF/DQykr0OLoyV78is
W4ZOLCnI/waiWpjXBrIByqJARaj4G93du9FY+08Dq8fR5lla0sQfSh+jIHo9rw/X
h95Wo6XfIEdmyOqYPxLRuSK5QTwKav/nyZiOEyhL6vOlC5cHwv5gxq1jP3M8s6OW
EOjswTf/ugRENfdPkouexY0XNQL1JCbDQFhyKi683Zuus7gEqFaI1GGXiHDWV0sX
r0dzGYcvzAM65H0tkKqUHCj8AZudKziSeW0DuJzbRTeMko/7OhoiD2V4zrQQZ29A
p3u1tJt83Rk/5lW6tmsa0ZMAwcj1tEMix9qQHZDJ4ewNj+ZAKGYOr7ph+G3PhRq8
HsAcY5Du4z9RA73XCBIiKL1amm073poa1+KBUOz3VEqlvFrHVNORERS5SNXqP5QB
9jZb4/cE1Qp3pSkIyt4JmWy/U/uBCm4R2aqEtZhmZ96wG2C5+LmrBxTBwm+a4EYv
KHcBsFxxlRqGA65nzsxE1cRBXosn+vb6l8xShOB0m4Ap+ee5uUD5GsaGMjeIL2Ip
DsThLxvzzFpBkbXvlNtLQGzNALfZ7hZ7hWVYF1s6e7asNALS6iN1zhv8RfG0wsgs
EpN9rHvvrcalTVkzFSv/FncHllssQvaMCyt/4fD2wRhZ006EFUoFMaY5g/lB6gj8
5yhty7rPS5IMKxupwLoEO3RunTOx1cTFpY8lr5LN1cNoa0QD0XviAMsfJkkX8B2H
gt+7LEgCiA403qDw7c40FAKGnhekRo7YoH75YFW71IWPydEazYs8BUDiknqabnzv
64E7Q7VkDdCPOcXXI8NMozBgsP0eJTBBmsr3F3w/zWyAsUXSm1oqFEsNDaQ1vy+e
arvRfr2uajF+6Fb3bajgknfTPqd0QHtwHMdBfy/qH+ah8voy/9PNMviCVVZpzmTh
9Ls5+W8rrUpLq3z0w5y2zthRvYFjLFsUEqm/JylPzFWLWkYQEHsIzE4l1JSJy3Hf
HPbAGcdkbi8jLEmZ2wnmcn8DA+APdWNmPBSn//fa1+gUCh0lLkwp7dnJ3S3ylcaJ
FJyvyHUhF0EhvCl4J9K4agijVBcV1GhaZICcev8uOfLP3PydcUcGI4QsuPQ+YgLo
eutRL/+rgMcbDmbgCVf6fXGd0opB0Pa+y56ZImHGE6RCQT0dWaH3/1QfdfKjrCM2
ZcMoDVresDV3xDq6mhbkOEYucF97HG+XzCgn1HBxNJcToj4jQ0EJypgSke6vg0fn
sG+ZitF+h8ws9Z5V7uEAoA6c6qJRE6GspvSZPzAQPwBht37G++PV6jK2C94VvF8X
brLd8fogyuDEU+u0ArFmCNL+8h8j2RR0b99qxIBqmR4sNtSFLnzGhXNm5mh+mZnk
bXDT7hVz4tezlvR+sizG2654B036QZW9GMr06HfxnjpcLWaBL45CPCdtbNEPfJjc
7aXHuY2b6QXX3rj3MBRZholPb0UDJpNGLibsi3Cc49ESsgNX7OShKj0NeiWQhugp
6OTrMrfUVaQ/XE6JI0VuHQpt7VulFAGE2x0faHJZvYiKUJYeVTKbeAdBD8s7Jw9E
2jei768t7pwEdfmbbieDXrHSnKbnHDW3IpEqE1PXtxaakvrmLry6pfuSPQ/YkPrT
jRGl6UN9E5DnfqFoL6EU97CEctvwImDAW9R9arUiiZUHNYDcmuvtVRnASUKQ9Yf3
JNcY8j1mCnXvicGvGu7pwYsK3YHdcDwuh8nXC7a0i6AuYQc6+k8izjzMvG2U7TSA
deJLyWZ0OzCXlj1ZqaARccDb4RjFiAT+N8VsoAmvbRcynEWVFZ+5eBaOAflu6nEE
9rDJ3eRgnc7s0nOS+KmzJFgK+9kN98gBzGK106uL5pyvfiuswei65NBbwI+VWTkx
MilEXDi9EQFykk44usNbphUzqxe8VOh8iQjYHadBvOxsNW/Bjd4nuRwIdS56c6uP
4IrjUNxNTKtSFoD0zQ0I9TaEhmtfeynWi7J8ejhHS81t9lQJAc9ZWi775CZnn9MN
F0gZobpdEhuxoJ0fn2dHJlOukDnvbi0gVWscLSBKgoZqA2U3lWKgcDkMK6+cWB4p
TjDeJZaTn0ByCxhCho+12ivBjOSs/86Po9kO6uy6pLN4tMJF6BuQJPuPr6J6JYtw
HAgJPM+q/LprTPuw4Z9nJm3/7SAfestKu5I66CZSToy9Emehgs7NQdyM9Du8f+ti
cwjOpvtg1J2F0Gc0AQfAubGUdp2wVlH5POUMNVdCjzQfMKXXd9x9g+QfUucGzT4i
EhXrwpe2XsylV2xHWiNVpoZWfXOjZqXBrbRguhoYuCtX/p1myEtA5apq4HKa0Ygp
ec7h/kLIDeiASAApNwshHvLOeNPz+lUKLtooHbse9qWMYOH2IJESMDi621kXrb1K
Ww3so7RfyDZhdhokuVwU0ITNon8fFype26fhRLk73ARLFXU80+/Z1AzX/ae1c0fB
JPB1kvf5dPihCR5/VtDWFBA1KEWsrfeiMY7UHd1UiaENDCvvW2Ct05rL7kCXkg8V
fP2k7S6pAJ08sbg9Vx43AXGzsO3Qo3yBMGx+wGtS8lMe0OxWYvyia3I0NKEN1/sQ
TJx8FjPfiAl+wvKvetA4Dq7jG0ParrfbvZmdNaBh8uflClurlIMjybDaF/pxjYt9
ru91NuFLDl0SW8y1a7oXBLUP30XyGoDw/m5Dd4z/o2ahIbUtTDMdClljjdwv4ZL2
QF/M1OePAjnXVNZqpXO+XbKbPeF0GcV/2RgKTx9pubpz02xog+sgGu8HLTY+iVDD
Pr/GFZ+Zv8R5bbE7EQsIL698l5dDErL9blOmPVROUDYskDpTbfXwTsk6ziwuWwhP
DY6FIFHhklMAoNTNfS3I1IG3dpojc/a+7jHozev6Q80x4V/FrUShQauAhXRXIu37
PwZBDIJWxaf4ffvZIP75PaxPrVhADWzYtN/pGUbUCSAtR+e0gNfB81sN86su4+lX
HCZzBWN2SceplHYGM9+aay7ML00TJ8yhsczn8juLeVii34Q1agcoCXUNmYqCJnpW
yTX7EfqgVqFTB0mrk3FPNxb5JocvVgwm+OZNKon4eJYDpO4KarGLMI1qsZIU39Wd
fdOQg3L1zeQMNNmwDDSCxZT/6TPJA3rJSTeqENCA4FPat8IJ25D4l5doPbp18yB/
PZBYxQ5j9RnaJXt2VXM0HFRZJopJ2fiITsiN8KmPFFakOYtgSyozBTxFQM2/gtZI
YcY6bCBo9PU8U+euOOGy5A6LYti/tLAzdo+G1u3QAx0BCk9zMqLBPbHZ1XzzHZsS
xrBlmLGoNmQbJGynCn261LZmSY7QlJsee/LOvZiCj5aoBvLgQet+8aAp2fUVN/c5
J5F7hLH+fyqyM0eTS8Wy7wRwEvUZ9E5TysQMchkz3Ko9HzSI8Ta7DhHFErhDEGHI
5LPP6fzCeICywGKd11c46SjhHY4gbMZferLTMgS6kucLlilcAheqyRQQZfwKVZkZ
rvAvAxCVigiMLverKz41CYrWIwiTiQWIbxYRWC6XFNVZNg/R+KcOTkbQB+rkmi/L
Nwv9g6o1oYEmkbAyeteWzUKVWHhkRRAV/bCTneu+wLc5t3yI0v8jagqAgic3tbTK
DXQUZFjd9644QEszyGpiSXDxPTA6okRksKZpXyZJw35iIeSFFIztgkm6qh1hI10W
CDVzpCNc553m1ucScUOi+vMvKBqTpK4E1YWL4CxRxY2LLuEQ/2MnnSDmZwTwxZNV
zQ1oRZDu7IERQRuue8Pm81BhGaIL81A+OhaMM48fEVnbiiXShPLhLTdBk8QlE7Er
JV4A01/yC7Q6YAQ7jP813dAFSJ2u+4ouhQ3AROiHASsHaYN9BsvHiMnhurqD8kt2
M/A70Ki32U57qq1Bv43k9xquVN+TygWyjHLO0yqaav60sUZdkOe8ZfpDpShR4ECB
WhCStXKWuE0YBoHkzO+pEIOe5vaDVJ3BKxINMtCDtFSjaf0bkmLk8M3ivvJILHug
CcExtGX/+1XMpFoDBDmQ+oTRDQkKHoSzDPdsOKRynN6Nl8o5PmfmjrGnio7VsQ3S
0pOS+9X0Zeqm5w+BVNF213zF4XU4pwkgRS8e4WCqy7lTkh8MIs+I3De2kehGbKCs
jW8qysOnzO9vMg1EKYEvwACoxvcwHKVgYl70dQGWSv2qyAizxjzF4zZNY2FZBBhM
wJ3NoZp+u4BB+Q2Usj1UgiXT1AYwDvHj4cKKdQFkLZJZvrgXF76Rsn0B85GodQif
1uXsQTdO+tERqGJ+MY56/56T/5N6q1GGWGTVWrHRSeNJBiuRtXjc9TZubNdKBbp7
shGnIHnNIfX0RvsyajNyzAOWFy9v4rsiufbPIUjBNoHBBSvZ5+2fsDhBLZ3/i3M2
zVDQgeAJ3AEshS3518rQIQnueELfFU4XQjcs0CdeiGuxVGET87nuCuXsf3zuxqso
giAO3MryqVei5+b/JussCZrce+iQzmo5GW5Nf6gLbYcGnwfsZchATBpJTRuZ5Pg8
W/p2erC4KFFOes00ajrVRwLFstdMWDhtYvwuBdF7YOttnIArIY1lcK0Ui7coApW2
TrkWtL4QEsDvMN3JgOen2WekCr1IwBR3oIrW7PApCa62mM2Y3ENjFJWc7CsZfEh2
rCvopRyq09GyliTwG6svbIyS0EY7bA93GsnSCVX05p93NV8Zhv6mQmBhH6aGOhs6
cWXpo9lGjQ67YhjeC+D4eIdroOsgVPtdz0YO2bHptB5BP9dcuofthlkZ+7J+V1yo
O0i3GFQVi6wc2Cwu2PXKf5acJv1pBHgiHVYgBac3bjNFzCybRT8crShyGd8Z980d
btQ9CISXIbPjnYDDfjncLq7xQRMNDh0BS+KuqomWC4ICgA6UUtCiD9fkZhS5fM42
Rl2HIXwrzlEYkTni2NUSX4pnCUCLkGbTZKBhCp8atUV3FPBd0WSoFb5pcKJUSbOc
AfaaWZ+sd/AJ+P162bsP80TsrvBGVmT7Q2Xcq7/pE5DZxdlbG6CK7cW4e1HoYl0Y
ewNo7eO3Ns31kuYfIysKHyiGMndX2T53vI+F8YE6MgtTlOFi/WByTnmoyJMUjj61
aJJjzxnaVBXCuR4fkPaZ+G4npw+7gC9iXrKUPXruBqQBCzZMI6+KUIoctcW28ygg
dVxqbqkqoEQJ29SbMBMMmHb9jmD2wftZ96vATwauv/AI1zXxzbic0w0oxzuJjqTq
8n4siyacvssMVlu0gDt2JexRLIzvHOFmp0tWf/1rItRRQKJKEdi2Y4BS9oJ4+n2Y
EQXHyvRqoAmPiu+0JAp6tC+zEqGg7ZAFuV3GN6fLzXhG85Zd9bque1d3SFoayqWD
HN+0KhVZDt88BM+VsgYip4t59KTCGcfQxwAInGSgQzA1pXc/PMqQqWB4A1cZLvT0
it8Wm5bFdgl+H++DrEJ7ptPerq53hnMST6HSFxSQxLTQXusd0xoqmnTHcwg+SeIX
xmHJfpcWZfJBjuVDNxj8CIx2Zwaq8MRyTofMOSHrNpH69AUBx7iosmK1fR/fMci5
uWQOv61MeIjdmIRbszHrgDHj+yepoIKYa50RsYlUSj9AgDn5UCFMUUhJISxySad6
TVvuEhOAh458s5qoZX+mxoP83Xh3+8j1KAWEt4nNRQQEdyanfkBO9SGC+CnZTOzA
TsiCh6pSdaurCwp7xLF7Q9uwxKfbuElJVTFL4JV99WR72bpE9WtTlvgocCukRz2L
K/QtPwFu8EFAGWyOV5oB+UC8tSUMZCk5m3EKuyRi+6up5cN/OpNVwXU6llsqoeWf
JI8027zcv909cCSQdiqHtSIyvekXbxiksxGDOCl5JPux2OQaGr2h1xzv/wFpWXxJ
P5Gr5nt0uIe79d8bjw87s/PtWuGdr2wteh+4nVVQ9OdxH8BNur8PmjJYtUyX0Zze
aR3r44u//X0+gANmMUFzzFvb7bV8YOZr5qfwLS91MiJbJ2Pbgcxk5m8zzRnFOtw8
acqPXFKMJpjz4gnqszBcONb/T8ridqFIYsBqM7TEahBqYrEr1dwxWCOIpfZcEcIU
rjCAViFrGA55MobZehpKuLCmbAA3ttytShsASYHLryaS4FVO54kfK2vkKpUedyxk
jfeNgIxslWTIjcWLXsT7VTHMHguZZm0NLmLwRASbvfJ+0LjhI1rJ9vWAxyg8nTFA
w7hE1TnXfU6X0SO4boKXI4IKSlC2+0nJyb7bOIwX06vQhvVLYWUYFinsyXNL6RJT
RvDH1DaiG9SFxKMnfNivglDoeT1MmNQ0UN76GupXHflvLTn9tk5O6gCoHNdvqzsI
OHxO+As2HSEyoX+bDoSgHpMUd8Tmz/U+nt08V2pAHfDWxzjKCyaz3N/ydjdt7Lyo
0r0YzQgo/5TOoa/WfJOdAD29RMo+6cnmmTDAml6LrgwjogkpYxBAWhMYOwHkYHPr
Niknel6vSfOreegy4NH43fdOqEkTZB+dOdlrwqCYrUiXesvZX85ALX8kJniZKWwu
TmGeFgWhYAqtfyhs6Oxc0jaA87P6sLcxo2mJ0K/cTkW1zJfIpmEZabJd9jFgk2eD
ZQphYD4gHZiyHsFqP+QE81JPg0BseL6JLluWUA6Jw7bp9PPbLFo0P6t1NN8db+aY
4Fb2YtTR458LjKnndNu0FknBTGxrTVi5wVJ3Ry7/8MIhE1Z+plN8vjZmfV8NWnyl
I17IDsWggxlyf/XrV2IHiOf4aPbr2NKYF7SNmDzQCSGKW0waZXqAzIaLDklzqg+G
nYLIuT01KEphVE9BrTJ63le94fa5Z5nb5esrLnDLIbAuHeiFlngexjN52Si+IiRM
ALilMKvNRY4/8P9Y7HGT2xnsVRUO49cW1slGvdhQaWChOQ8eeKp/nxBcA55nsvK7
pPYwgpdLaVRoybSu3yOsXAXgANLlcBUIBaXbOJU2NduoL/RdEwzTHxMzaEVEpVuu
bE/cvr79P31LdhwoO5nM9VOAPb1EhAbmmmfVBDSleXzLtUZxQIbGHgAqptIJRv4B
zvrgyRvaeFb9yFMTy0J7RvrsynWDJOBERv1XlpbKdkUnUGWAbuVTEYf+iyx7uhLQ
8j47f61Lm0P3zg+u7Rc4xxa6N3/Rm31vSzzPs+gj0E0vIrmL+pFVXnc+D/IXZPgD
ePWPmM8TunjFuKp6LScnV/CSQ7PYmGSw//gFe+s4Q44jUNiOAP6pT2xlMVe5ZUlw
847lC31qu4lwdZbYYC0jx5JZQ9/UhvYfRr86k9Z3z9dcbbii4ekazQLKMST7oH1v
eV8Ipmji4L3SaVpoRwhy9RpVz6ULgYXuCulAkOzEWoYd4VHBUU0OpFAkD0jGhoar
RASeHh40ElaD4uj5tqp+9QJ3eqHpiecn5ejExxAnrfe8TnOk5LwXnqDh2l7sCIGs
6N4qgu61glhHEEMS2ogER94orgQdHzqLBIaV3Tem18Qn10taLlo1i8VbVK+v/Cly
ypLuhtfGs/8RURmuH2oGWAuSW5ZpcSkd9JhKbhLSTtypX10tTjMtzzyCAR73A2f0
J7TatZtgpH9+HEycjSdWnGOFWrgeQ4MWm2KwjGESocLddmwD8qGqzszqbsQmtoth
wSizUBmjUOmmZH+f0RCiJQ==
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
OT9d2libKuIjCjBEvDA7fg7XeZek1nyP9hzlCHcB6TjKnhYMZF/9XdqhNqQ7PII1
wmPM3MZJibwhR0mOn0oLxBN72wmtMfcdn9b7Ze4ICAXzWivkue2VGy4TLU+EsGz5
hkTnFml9rCMM9zxktY05TL4+pvCJw8We8eCu8L9fBM4h/FkZSMSpx5GbOeUDRzGE
QJea6v+GfhXA7iNhP8RO6/6f9e030Vp7Eo+B+o8kj9Uh/e38HW2VucA8Zh0s5vTM
M5YdLMaP4mtz/BEHmjutKDPBRxPVUbGX204gGE+LSPT3D/T1+ALfInAqNlZsW+Y4
2+oZwNQW9hxIl5Dcl6L2Tw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 544 )
`pragma protect data_block
aAxB9K7H4vtVJUCIsVRXflwGHTldyUhhiCG4O9fYxbf3GSvA5ii7uGj9CFFvA0HW
OSEUR7CbQslC/eT1BhcORmvu3bnYtxDMLSADVJ9/EMe8E7PIy0KupKBJ8L8tYI1D
09+OYohN+//S0Ld8w0wyy3sbNwl/hlGpw6H1pFugXOji3klLBWjjzmmVgLcTaAuP
5SOpzGOI/YcAx6FUyXEVtzWtXF5M2BKhLsjyTjdcFlWZBWzTV/dlgSPXblVJ/Edl
JfwYWwjTunZmvZtLMi3Fnv9SCQn4RrAhv/B8AlGmBPp48wx7/0Q7qmjyRprF/xdf
4e7/uAYsrkh5MJFucYNd6/ckB6o+Sd+y9ckeaEtAujEcZvGxNFfCJwr3AXxNThPR
6F4SiOzFWWxGxi6bLrM6Fk491iDfBJT2FA2J7W+9ai+4kumsTjyB7NigClrRleXV
L1s2Nc4z3T150uwqsxOcLQKLB4+qqBxDsLjjoTs+UANhY4HLYBTdJbkn1pZ0WY1D
0zIjnHJy5hOKFiG4cRE0l+yTF1pCHBbepYfSZp8GYIAA6wiBuM+yk1dizALgrDC/
CkhsY6CtluKsNFD2Zq7H3dQuaYmhQVH/ffLs0D6nNJ7fwWV6RDiJhDjyWSzaCE5z
hJAU7sUuaqSuvMjIsptq1qRU9GMgZVKajLwaHgtRjreA+jsUYGC7X0/TULew0FKP
w8z/p3ExZH8GsYOuD82Nsw==
`pragma protect end_protected

//pragma protect end
`resetall
`timescale 1ns/1ps
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
ASlWjTZX06zJH5wZstUjKlIGBpYGNGHV3+x+sW0GeIYLwQKiD4xl06jjeBqjgxCg
RyrKWOa/qvTkJF24YrRqIvItjYuU0t1Yn3KGeftFRtS0TE/AosYnaC3Av6Ryj/+N
7rz1TpUrCp+oXaxBrxioGTUg066saVJWiXDbM/m9ZL+fhR7KzENAalgsAtzV+myT
MAkHHxIeqc6IQmFegSQzDLzYWsXUPh+nEaxCm24lXvmy6ll4Vrk+lVRGie1lstUB
3ax0jiQsqpktn0KRlsxBK6d834IcE50Bwq67b8UXDvHrbvONrixuetBVZhioNuH6
YDwQi+xY6glb3HY4ZtNQPQ==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 704 )
`pragma protect data_block
FnTLcw4M+YArQcEqw9HTUvCYgwzDSN/z4MnS71VC5zyMOqf5b7yD9DY4soouMfZT
HeJS0EFr/UrTDsrEuCEHFJWdfVmW5LraKVHlVeKrG0Tt0TV/MG6jxAdgvuS3NZlJ
rC86YSlPTUAshCBYeEnyg1IityGxKRWRr42gDR3+6VyfPVSq5HBAtq0tLBYnWJGG
8uorF7jYtxKm4Hg9Eov4LQubyaOXlwoZQD2gc7SIGVNL32eHFX4FC1v/b86ZsuyD
R2DUq4zBqWVGbRJGvfHLszLi6whyizQrIDkaWdxYmjNiJKAE3mL/oYOn7LPSV4sI
7RMGN3ylFIc939+Q+c1vM34tereMl17l0lHK3a/npli443A8TU49o28o4rJQSqiw
nPPYswMG3wyieC7yM2/m0497iJWguBPGxNOWFemwGsz36N8xzP0SXRwn+rvLj6rE
fEnkDuv9x/0l8jzEdKn9LYru9+sO8pt620m353hRMZUEfclSjiDhc9MbZL9IP8Hx
TVicdd5UGPnDfCgSP9zmfBhSKoR2Kn8EUXDrmnFgWoJZXvD1SvvBaCsp2CNh6D16
FzLjOD7LYYtAhpo1+5Tog8LhLDUBE6Ro7LZzkGmQpCXm+0ULG5UiBqPMsEn76jfz
P7FbZKybom8MnEadnMonud1a/6Fp3hlZWTc3lfHUL/Tp/6cP4fAlVbnEjk6a5kGZ
EJJ8ljFXhpuAJS3M/obitnhbtwkcZvh8VmtOrHDZS2FT2pERHfUMJfadU1V+xqPW
4Jg1+jZv5xin18p0jfkKB4zpTCOa5SMdIKbaNpjuFgnbvXlUe462CPK9rf5CQvfH
KJ5HnPR6JHVfkU3zF4TwjKgG1C/csgmWFlpSXz+aSw5KZAYHnvDCtEijlzRB3Bfb
mTZ8qz9AvORwspnFgFc5rLxrEjaoY+fuMjotsRp/wmg=
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
c5RogytI/ODELdpyESbtxlcc9J7/3u2HcKBsUSr8yiVVqKZe5Y2lzLQK6K6mshpb
MszTmqX4NNW3+77EK/2lK+rpAAp10D6vlAiVwOMkBdLxgX9XCr9Q+vyC2BmUfWWd
ta1wQ65DNB7dePS71WxSVHIqfd7rddPc+VKH1i2IYPJclDlhcw181OdBOIqoG6qX
F5VvVWJQjQCBe5iGmgvgEa2frmckscU1Y6Iohiu6UwY7QeqqOaSVgf4fn5K1S4TA
yDxqijPni4uXuKq4MekbgTW7FLaGx32Vp15kr7Yjc5XTUmSEt6uTfS28mMdRPv33
4g9KbiFIQdu4AjN8G9mQrA==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 7200 )
`pragma protect data_block
FOJ4tgHBCS5/epBsO/cA93qeT5TlfWhRFGMe4A5PkdONPzV8Dgt3ZYjCY/CoyiBu
D2gjbCcuVgIeO7B0Sqn+v/BsMW/GCqPet9iE92dVKNuR8pldxlBOBHa6hW2YobOe
uQvUf5hM1++x3HlgRcbDS+4eE+GUbgi3/WYa4PE08sZm2UIP5zgJXJUaBn5R1bOE
YfBPjOdn4T68RaIFcCTeitdiFbzrj6sKv821wpmF2VranTcUiN0v2jIKqVUmAR7l
q25nJ++obC9NPYjyZYzxUBejzNhHzvL+uJ1z2T9KrDP3HSt9nMTfUrbPWvMD3pnL
rV0yr9HykNgFCLXTMeRg9fMrSVjh6aIj6yHwlFALvpoiT1NlQdL8yKmrt3wb14nC
b8URDMWHfHWPojG1kj2amHeOQVOLuA/4ySAkDZM+ci1ZW9WNrMs65f/eykzEuMDm
fsNldlfYMuAlpAx38nzGx/4h9w5rh5Z00Dn6VRC8WcKWLF+rIJaSdH+0vjHfdQ7F
Cruhb1BDgcZCz+elGGpOiMB+2LCM+dAd/R8WVnILT+FS9Y7KTQpyu1yGthIeE6qB
iNrj7BbTjJ2n+uEJAeqJ0sAb9o5rA8euUXf/nX+AW6joIDXm/UsWHTPsbBbKIiMG
k8hSCOpFTXEWnqR829pqCHUkRz9ACGKV0ZV/aDCHZqKT8TTCYGizZQ2hxEjSH03C
BN2pNIhAe2xkqJfLleOUXTDoqVtSSP6gYqbSC+kKlVOrJdQhciG73ih55EdYoAF+
HzCFJ8m2KOSbG+C7Rc/d9Qe0KGrnOLCVEXibAA80LIyugLZDWSzXOH2fm6BjF0e/
ExlvCn463kfZMqL+GFFFJUknFLZVd5tuzRj4dWzbw4taokX63FvbA3/4+T+3LVl1
Ro8pOC+yOxSFqUEVPYUeaDVthc/qHy22pV8zpEbrSdEJfSmvLNZoen6aPvrzyuu5
IUBIzRYi82/leemO/F/hb8Zj8PFj9E8b6z+SwzjkPO+7baoDB0u7xliBPmjt2Smp
Gccpu0EKn1g1iN6ghzh5r4qrKMga6+H1Vs8dOfQLROdkb7rSSb/k4FRV9V5irUuc
+tOW7L5NK4O7Nsk9w9md3yC/o5akp1T1jBkGY6EYokr0bD7fwQ8VBmXxrStYWmzV
iQc0dYrxe0chV3L2SAXlFaN8DYO68c1N54s05EFR9Oviyu98lk5Vn6u7Lt4lH5I9
aVEVQOs8kcBFrAmeUxj8TkZ5e/TCbUyudTZXCivJeEySlJBhpsDqotq2sypFpDTw
bDk4ji9ApL0uGgN2mkV4C2BBwhThNPuEdN6JrqcEC5IXl/3S9ZpnHNmiaQLWczm2
M27yWQdmOMKEyueAnkF91h2R8u+O3X09jKtUJNk/SvXocOdBfEzW0+yxaZGno/ba
4gLJdDh3hXNaxX9KeXgPkJgpOV34zaac1RPrANuPso6JiBpsW2L36Bc1LmImkD1C
hKQzTiMSUbRul8Fw6QX7m06q4QtIsEqNP4c5rlRrECD5G00ac4H0hspV89yKKvsm
wceQizyb1YKK1/VFv/49rmWOjoU8PEIZsFrUD/sG7HDfDUq+1VwUUe1H1jaXVoIo
g6Qn6RceZQN7hjN7tFewXNL8kY20cbm8bY7CAC0hMRWMJqJ4B9XFK43iSYEdgnJg
azK1tLMX+MJqCmzwDB1imbLpEAcDSxsiFuIZyAj8rDZxzxlyqYl2um7Kh+UH8Z6r
LnkflLawDs/NX7DPtEZrO76ixP1kILIxpNBZUiRHB+j3g+wKx1VFPgHkqDmlq5kc
M/4flHVqS0L+QPcXvMK7VWQ9w7uzV6WTK44NGBYhNowTqXaP5VZobU64BebqaOUf
oRLlz3upzDe7ZXMiEkRyXfiXmAYa3JKpfnQR/lxDAOndie1ewezhtW/OO8plYFEl
Zr3ZDAMP8Wg4pIjM/NvoRGZYKYNy0IbGaGniw66CRZdjvFWW+ULhsbWC/tNAK3nH
tHzZmgGttZJ8dhEZ/JF2yaI0vB7qqml+EuMfUPKAJv8zFk+pyOA4EpF/oygrO/Bs
tscG8HiR6cGdz0LzGw8c2CRuUiFNpjryWgRPjsjig+j8OlB3lF+86+4iOTJHQfFg
P84QybspS+E8agPYeGpSG5HW6kT/lM07IZAtAoMZKc/nMB7C6NxgwOVSX5vmIbMI
A1SWMRXB7IEyo5pSsJLZ6W+uCDla6VDGIpsyyCwUPyQqDyLqKM2SS9K85IGRie4u
3y36sNf2z9ZGhJ/xHdaRecL0rWOpObE4KYpuHNr43ipQN1btwCIMgJPb+NTCvf4x
KgT+pBBAzbcvHQ80suZFDx/hV8VGeUTwPqjL+8pBq4BAavQB9/6//6pbRGzY41LQ
38EhcdR7dgbqa9c8rRBi1h80yucZilJGNO2ZImHANVJlL7dFhhNWRvKaBkbFVCrd
Npvn0LrGhyn4ggbQa+FwMQZ4cZoQGtxrFCvURfgxPlrW8yJr7G/94+9E/EUHKptn
6LatEyyMPYvgv1u4d57JAEZ48y7bSsD9WeKNdyMb6+wsiefplrBcMki/XE8F3ROF
hD6NSyJzO5tcMc1QsSE8XY9gw0V0IlNGjuc4Xsj+VfpxGJ4nrxoFcV6iUGzFR2Lu
K5wFV1Hk7ntinv+HWTg2Rjl7zbvEZiGcM9rdcQCESqY63bvfUVy4UHYi0o4Lig7k
PWV6lUVQkIK+mczcXfHAdAi7sBdEPsC+tQANhfhmqEqshak6bZGTuuzKmUgBKZ8y
hiqEPF/3cK21OBudAC7FbeV/0nfsLS6AV4edhCdt9iYjt1RLh1us1MrzO8nGwfkV
LYmE3wZCs+vO44RqwYSXHGl0KEl4v9rheVAd8Uvqd1aoU9QXdiq+F9kfodW6eJDt
bZvaqZQMVpdmIi6MPoL8oNkGWv3Sju1+rvHW/YbAtgsCCQtCeq/+0KZ9OTJaeKvK
ROuLoUD1ec6xaWb0dmBPX/fWtOS8ojSLmdCx0CPWgoAEmI88vWrlUuEE5hfy1D2j
SXRgzmymdn8ELUGfKKcOGvMFOCgFhNC1T+B9xf9/6rMxxG30YtlyCc+cE71jITRh
fY0Ip5mH1YjkjjtFHK4WYj7psd8zt35zsYIYHlX97xyc5PF47jQy8hIZw7dl/+zb
OKpQt6aoJiDhZfhfEk0M49Mbmd1HNRuO7OnqlA87PzTLnuGZl7v8SZOrwf1alcOl
65+fkP1lP+quv070PGAs6dQbaZ0eHu0nuI4fthJNwUEG0jo6jjz897XtX/f58d0Y
iUFV1aZwcx7OlrsA2+SfW9lHHTIIear4AjT10PzjDlcWuYaPlwE0U7AdDAqQefLT
NGI7x3izfdaLJL03CPH2MWIb1kF8/BwtXY4yX7UOdEZTKOF5H76Uerh2ZBYzG/2x
hnxds3ZffeJEpucFX9NPIe+kCH+ksh6cVPCwj/A2iXzgqSBvFqR4aBkjfVXpAhiV
lDyL0LOErvGkLDbWcvAsv4oZwvKoT/oIUJ/5Utlq1ie+R3sIQDmhilbQE0RV6UbC
gZCMyDwzg7RhrZsJo1H64Z9srG7NgMxZXrqZ5ubGbAIEpTnrxqD/XtnfEZ2Lu205
JSIdcB9W2dxg4w9xRcQdN9Oexz4YzfRU8FP396pb5UZh1y/w9gaIfkQuy8d79gmG
2PnMk8tuPaTFg9UGI2E9Zwn4JiWJ440f3O56WtE/brI8f4Fc5YmzQOTeWYncVB/s
G95b6q58nxM7geRGCEBZZKc6MIQ4oHhuXlK+E80Kij/1ffSl2rEem13nAGN95nf+
BPZ4UqxjXofIpilJAHiUNziGG8hMP6el5dDRzNgHDEEzenq0CH8E7KjU8wgMfVJA
wNmqMRPs4qcpsaT+fcZ1JBrCGcCyqq5DpqJEcUf6cWrgvuzETWmOcrcuK/q1K549
xZKUfhYBKG9I4sGoKZmQf+PneM4IWLO/rhEygrsAL0gRkKpmBOSTa9+N5W75nPzJ
PEiQNY0iPvYnTdTS4LtD82pmH+5KUD+s9k+hoCtN3eNHlANgf51lUXMFQAkSEHmG
GyENC/XN1f9756zmQLlDUcsfIML/UDYbYeJr1JME/ODOPln/tC44M+MINeJbD6ey
AnyWY4eZxBoyPDtu0xeS11UN1gwdR+doWUx47Obml5zCJFYuifmKZRYW+GYfWNIR
QvBAyaEW4yhvUZES/dN+UYi7mJ3BTGbOmjAjQkeFhTDoaK2lfq73h7zyeAvPMtvM
D5CZhYtAdpcBplT2pLz3e/sOrfexpgvZH3CNI2GVewGPf8DfzDDU2dPuvKfoDKls
I3V9L/GUdPZ26hCCscsyFYIqRjXxQilC4mNB61oQosc8lsFaDJIu24+KVocMhR/6
AFcY1b67xzmT5YX9aom0sCYdQcqeHaKxDliXrL7WgszlEcHfd9uLMC5Ct+V/dKps
LvuKwVa2D4lF76QTrTfzVEFufYsDZxo0o9ol1En0KoFQZkxoZQn8uXv1eni5T+C/
aiYf5BuL9yPC5qyrqYIYpRckN5TFRDESfEhceTjDbpJrqo0uiH4U7zKmkL1DA5av
SFXvKAApQxVuJPnloyPIqq2IocYUm+q/5Q2o67T2c/vqTe3gbXhAT/AAEUUJbD75
II+54ov3c1kHT8eKi5vonWMIP9Y9EidY1i1YKL28dutytLcwi6rrLesT967aysli
x1kIOiZ3gvowJ5YQP9aG+T78WaI+vUjWo6u8InrtAESSzlkDoJ7L/0Mi+oreoWmD
jUgzZH8oUqcG3h1McFPoEbMsmEPltvF9zKbmlFPtEvSWuZye6v/+Yt5k0F2Bx0oT
SJJ6EzMP6kt/C3LTyu39dQ+dm04TSW0CnEcRt4r5h9TSKFGATJ2RYIT3GTVpuuoc
Zx9xy3rlLcbHxuKFj4L/KMQqre/XO+SpYp7R5QiOdeTMQeO2cil+xZXSUh5/84Tz
uLaXj4oOjrDfR1gbKbvGFC6N5OownOfBEI97SaZF0t3ojchqhUjRW3/ZIyEzbXze
/YuEuqR7LBHcVVE9KbexjKjpKKtACVws1avPyhnQlbsmVTbD4ISDtOQAFLHO3EaC
59vwQvNPYijFaey6SY0adiDdqmg6CvQPEhWyHa13HvRjXt1t41TEMJsjPDnBoG16
AvqtOxfqIbKIn3pzrLhzGwEhw6k2XJPpI7HDQs58r8hJYI3DIfVjSzBv4NncaBlh
YzAc/aCS6GP+K7KYKGHUAZh/BU9WsmlkI83rlfioWphcDU3EsGJEeFGBczs/ZzO6
rZ1UE1Yp3y57qIUptYtxyy/jMcpegm+ljtoYFnA4CVpbfZBRutDjdJcUamhiJFwV
ofpSp6AjFfuCYqHWOOcOYJIIwMPbD2Y+aUDdWUYqZ4KE8KJW/P9b5iKVDth2ax+t
m3yEjYGJ1//6RDoVZgz7SfTsI4yJSCBjxTd9YVc51Ej9ZWoXr+sd7jTEFRKyN6v7
GEOFEW5EX3v+Lx3AoD8HU0CrL2xB9TzV2h61p8mBZ/8ufQnEDTNrAXOaqXr3Ovz3
hcp/Ht+nbxzTxjqoNTFPHe2Z6IZOKoLp1Hzh4NA9pceFCs+Ym0K0qh/c0Yh8xG3t
8QhBlZVyTbOB+eFPMf1tftuBws5/I5MKqGq2aANfT9SOGjfh9wNNDlS8CpH8ZGpZ
NX/MZzCf4qR6Ia0+YyGalGAvVRUtffzhPhkkrWsQco5tvdmDxRWE8TWGpXu4zzPz
7NG0V3yMXkSHXNpktyeKVVbY2KC3j/9xouTAWQFX0AdgXxecubYE2HGOgJCtgWHA
CEmXQpzwu1zXutOyyKz/GdtlduuQX6GvpOmD0d3Yw2sL15zcLYzPEiZrwxO1W10B
WnS8qhoayfji+Dx2Xc6Y/eDITCzwf2xftRaI8gnCBT72QcnxgD0vM67RwQ8UPiWp
yiufgmc59n3pdTA4VpwJQdsKJpuBTU5jIvAoiLlwheMNnJTCQ0jgXfEq4ZqIzgHF
e8u7YHYU07pnDj61AMM31UuTESeTefQG/GEXlggcQjcODoLyB7noSpl+jJIox+Cj
Bq1lsKXwGe2m+oDHThAz437qdTBXi896yXwXjjyu9LYawT6kLfKRFsZB2kw5RQK7
VBiQJbd8zUMmd9TmJEiCKJOcRylRedVNng/Jk4ZsxtLiYX32HgMZtOWXFgZEb08k
rqaC8Islqx07Rd+JhRdIAGVz2itx1+fs+LoTbrrsugSi7qMuyJwfVVoChPqzv0ry
Ol7oVtE2IagSz/vCA926qcOp3KhnPUIFa30rAGJMn14Pfvu6FEn3zSLxVp54l9Mk
/k02+w2BJklYPCECW3rkpKigZVnOwomFGNW7IxjAeTV9J2Qiwwiao2zU6M/bNEas
f2rdRYPp1SS3ImHMUue1fvPdKiwzpKQq0X2rqSRRHO8AjlD9pzwVg6KtMCBBC9l4
YrGd/z2DIN/+LKesBXYEB5F8LORcMlDlBpWj2fSc/sSXM6+q9pdiDd+8JZdN7+uK
DnMmwNw/8l4unks83mRXKwfmUee6g0Od8D36StMcZo2CHTtYBsjX3aZC5qwJnunS
eZ2ilpPAhRdJmr74zOQakj1sncSiJOz77v/2B7VxFzTim2ih6V8/dPMXOMvMEkeZ
VmJ+5jNbIMsIuqUJUfHH9YF1nzXisISZEEfosIq0sB7WDmQ4yHRCSsVwS9BFMbLD
Vps5JChP7NxFBneGjI45iIRzuJfikpXT7g132QudC611YA02vY7xSxH6K80Ev6a+
s0an5GGkoBEhAby6FerQL0ast4DimCx0IWaXleMizrgYDCl6bmq8glvSHrweznTv
60cN92lbgQLz2BiTG1Qdg34O/HEESg0koRB+93yHhemzau8zrMuYMasvsx5LGQZd
yo+TGrefMJuRnlt7DGo6ohJW4FSb+H+PmJHOLs861ZnArscFYMqQnzRdU6pBdtFT
Fx1zmaJXG3GW1WpzDUAWKf5883VrQSioPstlSQ93XWoGlSZjxpNWv4m8ofJqGPSr
PZaByA+FgzYTeqI1GNQT1wYfC7HJAawy4LdwM4+BHlAM+XH2IXCiCkkjl1iKb+BF
0MycLnhdT1SlYuuX2Iy+UN540a8Ory8vtEDLrH1nJxEePQqnZmcfjZnE2EQQtOpm
W61ySV3jrwblsrw/pgVrGoN+zhaQmRZLnWCFdsEsS6PlidVulTCfAK4xL7zjhH0E
vg5eyamR6brdrQlKsSDQWYWZ85hljjnMkuE3eKg9/+/Ia/8e7kEsLHgIi9+/AE+C
XrLLgyBhfsc2u8AxwXVFLiqcFNyAoNHrcUKtTlejoTnBTBGOgFJdawVanYDEFS16
+0l05IpQEOniS2MqsiDrMvn79fL0eRqFWY7UvmfgZ8hFPqZWTZdpIbjjQcO+/4U8
CREZcbPIC5U6b0/G0xcnN5YF17dcjqXj3/8VBdQ3gsZjSPLe+J3fbNO29OCrOAyK
Bc5XH5YdFlBIEME2y/gmbQ9fpb+XVDwzIStBbtAaIvSemY/23+ts7uOyhEGDQBjI
+uKEZDJWPXk2c0iYuGGkUJSUATO1MCwiPTI+IoJu2TcDtHOJRxhKFFxf1XOGrcDG
hPKeeXijl15zUlBsyvjZwuCakROO169HDocGEqv7S4FvcQbZVjzj13dQ1yMLfkG1
sIph1o0FIJ2DbZ6GqA33SGOvpUgsPno0NSqGLoRYwhTV3KMLuT3OC7bx2rZXf9SO
RimMgg7/mVOqvLs5ZTdejkneJeX/xFlJWFhWX4wdyUyE0/07nKIom74De6LSJCez
9yo3r2nY3ukXQjq0PLVQwjzPgVAwxBSfNGvcd/woBQqD29w7EzIgDtN/qLgbqRHP
6hEKjgmNsa7p1m3OwdJpeYr6CvNePWAdODyBBLbhAGP2y6PfA2Jk2SlOHA9S38bd
w6iL2385mhyDXCqqEnxULoS/9GvlD4WD18PlMLIfdFxNxpam8fK+TFINMHNsHLGC
rb8sGLjeUjCaV+U4Kdyv2cpSTukWJAdzqCMFBR2loSzxsoAKhkHth8lYPE1lq4TY
Ja4WaO6WpJ5rTEz3ZCW6PnPCI4sm1p1OgutGImo+volGWfQZCoGZP55QbB3dcryx
OsC//sZe4lPlr7ewEbLJvCVFbUoxUPfAF+wTJR9ArxmwLEgCz6Qzgrw1wPPDGbxe
Z1L5NAP1oktBq0Md3r4omo+0/GxHc7AFP+y0QNRJmayAnCErZrnXSE7BiFtZCtcx
UEbCeHYx0YGHaDhzsHzyiCve+g+BKaduTDh0pKuWRoTzFnQ/Jurjd8UOcRQ6W/C4
gVdH1YZSw5d+pcMOXdIPrBpyg0aeh25wyXddeSciLkaQ2bFVAn/KgJ1KJUGqM22j
RxSSM/asEL4A8Ha4ZOvzkNoYOoA++4mm0JpJz/sv3qV2HGlcVrJNCqapWXrGjiyr
pv86dbnwJErqYEdQS0B2lvZp81eE2s2+FPNABNowxDcWbXnXc13SXjMDQaO47Baz
s7TR/Z/hIoWp0U3+0e7EDg7i+vRM7WaaMWcEE2ovIb63bNAMQFHIiyEpuSLusCs2
KBlTo7/tD0lk87cZWY2BYlBitLCR6j6YhvGR6FEjSyQteF/y+RfwY1yyVsUJIhhM
zIYuyu/o5jhwnhFpFKnS23nLepvrQ+28AgK49fcYxun57sd9Oo+rHHVGdNoiXuCn
B3E7NYe7E/VNgB4HD1+8rO0U/iBnunncfhs3rn908Ca3vMRtIeZT6M1MSeo9ipbO
jN7PvG7bgiYufF3ZZ4FmsGf3nbyl2EMB4a2tqhgHD2E8ZgIGZRLa2IIHzLT0k9Sq
pWmxGE3DbykmqxGp+e9JQeE0oHAQMWAdDeOwdfXY3/V8uWSEVwfscXu0bweCTMtB
lGoKrLEhnvmHS7O93dd2zgyOjqQVUR08G6K2mei9BUAmOlyKjLQNRkbnnFqwlGV9
3w73UxivKJ7hB1/4IA8GPkjWW9wSgoi7YRpHaQ98tL1vY42bI7etU8pXYhWbeTYQ
EF1dLY82hCaMoZZJP03zeNddrPbrYIAhS7E1vgOKKFhlRLWmjVWpWIMBAOemzgXA
vwEGA+ahx3JlibySRAULOLUUjcfDQS9Ule7bGx12pwddovjisGPfWVz4KBvmXos0
VfRirYKQ/AwFelauSsbdWmoTIKZkYiZZuefmFVAJKvEJDiBjXH2yWUpyNJ1zJ+Jk
21zJIPUrKgMJC/TS6U6NXNFOAaxpTOA4Ff2R3hhMAqmddUTGgKfQ7xQiYmYmCeor
IGfZGlQxdyTy1KxFehv3I2B4QDy5DF+gfpA1j9ZL2KrQGteQB7Yse5A+hKVBxZ0m
4hm7Q/Ndc9DCTKF7gPZaDfgRvCjsCKi906ngNzMN9VtjFqYCrOwgzLYdBmK92FmI
9NGV8R4Q8cYw3WojEODnaBaD7XXMBOWvlbUUtiVAKe5/feKHk4gBxp9hr0F2yPzo
VENEE/MNeCMAj6ZNx7K4BXe/qu9rapC9b0dsWiFpJK4k7+ElQcJYIMMsZ3zJ7bey
rsacLcnpcC3xO8Iiky6CSc7mudkPbfDd0DHhiX4THIs8Jngrnt7kRnrfxWLCpJmc
jdiKxT8oy3Ahz0D5RYYlvQJGmb4rUhxqQnff7w31vUB+n1Gu0Ckm0yCirLzDrUQy
`pragma protect end_protected

//pragma protect end
//pragma protect
//pragma protect begin

/* Encryption Envelope */

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2021.1"
`pragma protect key_keyowner = "Efinix Inc." , key_keyname = "EFX_K01"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
aj98+imdCHgwEiHhgsXb7o0EdQLkk6kgT0V7mPnFbv/sj07MKSCTAfO4811Kq8Dv
iTMypygrTBNbG6iiAQSIKDcnw4gxt7s7naHRmfaLvAo8O8/2ilH8o2gOmVLpVda+
cEsNEmLeiDqZpMRUZWRhNbbM2OTfLaHjCHF0ajZxgw5A9kBBZUcfqD43Xtucd2ND
+IejFeM8sxitLV6cmLPFIE7h7PQtDzoR2lvl6OINtgPxn8NCM9pJIbBcSjPn7gQ7
TXHTf6rEbmSup7Dz+hoytxrDy2wma3/ZQG8T9sd/NQn0YzUjtlKQXcy/D+YQbo1i
GsZ+xLDLd7D2Le3IQkiNlw==
`pragma protect data_method = "aes256-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 9296 )
`pragma protect data_block
uYj+qiom2boC2X+aIjOyy1s+DVXysyizk4pVWEQfNzLfPxFXB1m6o6f3Hpwadrix
YJw1Gg5q5maAMH4hY2GxGMUcJ9HRfsRmKopEmCsilS1vWBD660QEXz6kCBcVhfFT
JNHyOzS3dMu1lt3DiAu3h157XK/u7Pz8RBAu29nRblJ2yempTC+z2XxFtyQ5BFgS
ODdkl8nsFx5CeQcpXmaNF44fKynDfM8mdkNbIU32tInsJlNeNdPH+vAKNRlsseuI
chqNTv0ib/TnVGymk/TZ5/gwSbINCBPFRRymxTPXNoy5K33fbtc+dLh8gePJh4cV
eKItzD9gTbcbNgfxW+bvDsCiuEfbnQuxfMUCKJ/jHNrAIoXPhvWjQQtZRKJa2mMY
qIzrEA1qsx4PL15dScmUIe610DCza5DDRKgAcqhl8rJhIWsOKIcgRAnKN+y2P50C
K0heK4jLZHW5DOkq+CLVQ/0q8Pz1TnmsWTPBhdmhQCgSsTQ3OdEH/toaRZn2Zo9X
eGvUz+AnAHyZLtDFkeIxoQ7pAEuRnWFkNOs8ANo9+usQ2lvFru02ao/P4mh+WjWP
WZGlROwjm1DCXxPQrkmGKSpJUnyiag0alD+La4EyhVkxacG3KG2Im5TPMawcrHZC
4Wn2/jCxFi1WxlL9NsmVSnS3vWm2uKWuMygLBuFM4PVgY914XsIUVxtZPfIokeVR
2+rDbya4IiEvhGolRXc52p2IiFGtZBgZpKwaH7ZXQYW9i08wvptC0Ax6lG+tmjRe
fJQ5lAUIQf3LzMKWDkH90Jc3B+lYkBCnnyxYOQu6jMSapA0GX4pdM7gzq64X++tk
YUg5stIK5YNraEyYaot6OT6+O02COFu46qiPLqj+lzyG3V/OAyqc1t6OBbht+9Fu
0lYhYK3kg0jBojnfIGtCqtIZTZnAt9ymvJPa/jvoa+bsK00nRLdWnYcVat9w4A6K
KziPgAjxUq4FanNe5kchdwKv8tzQ2mrnCJkPWJQcMgYf30VARYqTzc2nfo+RtpVG
QzHnxUFZTe8MXymiHBynSKxkyict/DY8nUBoX2tnzCs7qdNrNGoN00M0y6iSggm8
LknOunrhsU4jvrxAQT5mz3Ih+4DwzmXrBE7TCVPXurTbxi9GKK5VmED3wxUQQYEI
Ha/aG07Aax4PUCE2bXRnVU21wGIg3hARDKVsVsZ+2JGG+uJHLmhi8535t1cn9z7O
Rsa7Ru0+o4s+mBiaL3CHp4lnQNINjolAwNApjC7tiZWAZAr5SB/uXHUrRTZuDFXA
WBnWYiZ5L2nOhkt9ZDTuPAEVkTF1qplMXa72k+O57UTE5NvrxtwzSfBpbjeenRGq
zJ5Ge1TFby8PtX3aIMq0JzChQU6Pa/1UA+TK4jl25TLka5mQawtaC/+6dPg7mXRV
TBSI5hUdJ5KvIu0rsFaLJav52ru43xfX+o+n3zN84P4QPDStBUl5tkgZ+5SBW4HA
qsGs8UxJ7UzQgersjOnIQtWXWxdl7Z/8gjCf2EqFWxfnUjrRqZFE8fpqFldI7lTq
Na7qvTXkuXZjZi0IjsQi6vxrQznH7g6hp6NMl7yC05Am2mVKTwRfHl58KQtB6ZqF
+4VfE+zA0twl8AKWyPy3QtN7c+ljWJu+Y0jJOYh+Cu5mta5m/Tudc/cShhCaBla2
qUXsjzdmb6aj99jyCuQ2ZKaIznctxQ25SD/cYXiwdGSJ2B7E2WYN3rmhP3Nz7fuS
BJQ91vIMjg9ZJeHzMJERy8CQZzlmszCTiKWkimnueVLLMEkFeQVB0h6iL0Z+XvzL
vhBFWcMhAE9wwV9hTdJaw5CoLvEjqxlAuVFd7NEcT+0WP/X0uBzZjxG55ZtiFPM3
6kSdduPK6yZfzrQ9hiL5YaAUh0fCMlpKgCwmhChbqKCAolbqL/vhMi5RD0Oml59E
22PNr7AG8jMgFwgulKap01RWgf34BWhZRBYH+syOn46ls7Oi1tDZ40xYxx0v+8UT
WJDBnXhITTJzk+TplcOhVRmUw6jLJXiLiyPapbID9lMI1jnEDEO4AZvDzxdrFZyO
k3qH0oIXnejpCfq+BiACSVqQ1o7Ss5ZE/GgFUCuJhJVCvEzkB8WxXfsLrCIr77aL
nutD02iHIbmb4uilsxnignpqagD5jEstsNJFimht30ZUznDKX/J8O97enpgy/2zi
KfWXYVZSbSgLWn5vrtj3NzR47OJejzXw9V7kXmKTDv9Sl6RK7mOXNWeTLlaOWbKW
GRzjPY19scHGOn3oPmHq35ymLuLCbD9sc6KHjYBmmgrV53XXMON77XCNMyiqC+Hr
deoHRgu0A9fkW7Ch4/A/9DwydGVF8c59iSzPtZuo7WnAqLrkkxUvGZsqG1pOPSpo
Jooq0lXT8Z1IyP29gceMsETUl+M4e8cqrlfvcLB5E62E/keoKoSJfbK43DoLIa1+
JlcCJJdvz0LPhW+vcTqWiJ/VMZCwUqD0+tbt1efzx7Jh5tKAdoZ54+PICw9ULs5o
KRCoKJck1yDqPCDrv5srxlX9N3E/xvgYCdZS1vz++o/SI1njPwxw+hjqfDN3gNHN
gsafpGEBMLtMC7anYCLTbDTCUeqJOkBmxelQK2zfpMU4zKfslHdscsiCF1CtB94c
xh243YbcR1xoM07vGxzYyFz7qAmAQQwpg75Nq070d7zCinWOczkDbsfTZfGd0eKW
WR30HwWUnYcDvNRCATzm1sSFAhA1MSW13mWQQR9H2Gfqqn6Ecwoeh8wZq98hYE2e
dGxiTJOvSZtekQjd7R4za+PLTh6GgcBqOYGz/kkcwLMQxBcnI72qZMY4K8eQk0xW
/fIne8/ENnEmbFAUqIa88pZtVay04fbV/4pPfoYL67KsTg2zGejSqxo+tyQdXtbB
IX7dR08yJFb0tI4CRrcfSslJHmGUO4o6PqPqI0wSegcmUKCO82Uq25IjwYxHBoE7
8ITyx0akqHq8F2BvOnueSCLIbhEBXRn7AWvUOxF9CMU6WPRmMH2UKfoMM/USBSp2
BS670U+2Njso5/pEFOc3ii4ZjdEk3UwOglaKr3/HTUDv2Yc8Y6Gu7LJnSYPuKbRk
JBjpGRFCwRrk5ydl7CU7ED+T7xKibctELSI8DRNanOgZ3l8tfUrUvfLHOfKNtw5W
z53Dul0TkJdQ12vES0YApCb+QridZmNiU6mT1k2eQmmeKNYIHBVFaiXXA0AmzHJ9
pzvM84vrGP45sDGZu2HFSSlPI21NqEDGbM44z4ACi09ojAnvrseNb2RUd6WCWUGA
mSo99e7xSlVeu4J1XYi9US9YugMcE6xmDZMeKrZOk5MVDVifeCDFU3AgzXhlIEff
J9BYwixWtrUZEPqW7h4rbzTthW6VBN5rpIaqjgKJD2I+EKhmk3AdXXHmm2Qb2P6D
lkxlXJ1S+v6kHlRfvjHdDTHeDUVxNfh1VabWG+x3LrP2Xpn/NjV4xNQQxRu23dG+
hU/K76ZSYCKYBlXlSpMWTXuchtlOjUn2AlHt1ESHZMHTzs0ljJzPLY01DzNUvz/S
izVsAZLqKuDkCsfP4YrD+ndyPb5SAXBl2EmanTqjIWaVaOdYSe8A5uwYD4qBo/eb
SCIjkb824M0u+3rZE8bJEOgZxyP+vTaGfdDDFyAM6fXdr2PpiAf6O41T9Vszc1EV
XYeDyTlWfASRm7fyL2W/nx9pUY/gxWFFBkBbNZhuNPwfCSaCEE+xmZOmpUsP26ni
ln8asr5H76nOJsZb9B2fCr5rKdQfIPXD7/4wuBUj+uweqEARYUyGGjP00MmUkv7h
Ikm1B5Hmoaavhrlt5hiaHZv6y4TN25fq7gIPglv335UoXOtSNl7VQjMXovhefOpL
EDaOA0M7FQj+c2wsU9fKNE7mPZ5dDpixlk6a5GPRqGHQRQZBRp4LFi2WZaBXR1jy
wlyWe3Je7iGP/8Uf4iee7VzKOVU3Q910mlqM1bMrwLJrs2LMfA40kfxfxbOsPVT0
rVgQACDS2p2gih7OMoWPTSWTndTHZ0Y4380O6g4NLw/0Nt9faxnHpKxbT15mCGd6
EL1yepl1mLcSYEoFwr4S0hwRCWpFHOgN4so2UzNYbCiMa0024blLjoo4QXHNYniY
0YW1VFQ2PcWo9u5ueDNdQrQuXksC5qv9wZ3zCCNF4HkKv7zus5lmJRYi7cF5yEDY
rkaLG7iA78MMFugF8TcV9WsIFOy4EaexAivR0jTTBt+UtE/QHmPL/lichA7SmaGz
wziSEQlHrbV0HS3F/7nrXa1D1m6d1CrBcgJaWIjiEJ+EwjPjA1VdmxxgrqHUmku2
VVyMD0sHfaMNmkhZC/u9E1hgK845Fn0FZfg6pccbmG95IioJ+7MLE8B0+nH5Hst6
UyelsPUap31Ym3pnrfQg56mXRJdFQSKdWhtj+y562WUnvyJAFYru/wy2v+JDdi3x
9Pb54vtDPjVFi0Xayq5BgwR0SRaWbWeWqLqHJZQmL7lsrWU9UQjHsX3IlW26Emju
PsuXXL/oezItn1sKfTLitlWHcqQeZ/6tWi0nO33uDAR199jj/VjHih10vKYByK6r
HHZ7+7uYZHPavbkEGgvemBVLF7+1R++smN+vXUk+YRWSGQnh1Th+ZVt2imrF/zXL
k9jjoW+fe52nSnvFGHizEeYJCs7RmilwmC/WUmZbAC+5Wcz4AXze+u5dc9ptlhM8
k04lleE+C9Gt1R5soEz9zRHkLn9QhfkR38x2nlQ90VnynG10bNRNNGXDCRe980DJ
+qqgCcAiwD3Watl1d1w0nciUSa36O9iFA+nCJTOvcOIwq/xJ9hdwimCkLOf4DSE8
6hmAoImb5AzH5Hv/yfoVcDlXzGD/5Q1lkApwb+isn+CkdE9z+jFu648mabhIw6l0
jXiL8EwApiBOX9F+YjNuNG4GifFGiTyAK2Bk02Nw9PyIdUOPuRzOBIZWCOG1f31g
oPaVUls4DAmcDPRHg9ZukeQeHRwu6+kFkEgi8VxMbVfXwyF4rfNjhnLq8K/LVt8w
8rsD1r3XVpnySconSN60Sa0eWsszy2Gnf93EWr0my6XpkOsohN4RZ+mZcrTZ8aM1
mKdWpMJxw+pvLLDNoXm91PPcBKo1xae3OUOYR93E+Au/U80Lx/D1Qn7NOSniAkUB
rNibM57XgYd0hf3fqGFRsTI+5cBAOtNscPVt+mSzG6t3Y5sbNILA0kUpQdQzou3R
MTKY3dm/H21ZAS9tU1LwM2xCaHLiqEfedilBom3IwlhBNJEqRkJv0CeAec0TezO0
5ZvgSQ3n7kKkNlfnWulGCqS5vpM6VLXal3WH2aRNBqDtjB1D/r0w925kWK7B40F8
eXcNthpSqoXq0mIA0UwsNr1DJyGDPqPmRTghZa7Ro7Y6MzXryQu8qQzlUcBlcsc7
FxeOiccQ2YJg6s8kM51wyrqj/UdVX1GvPIOGgBPPD6yN/6ABc6+7LE3C5z2lOKuc
kSHB9GtS1Rpa+BTjp83lFnYoz3x2WOm6H+sAvtbEZfHEDro/Rb6yK6U7MEXHoSRE
hLWMGpMwSOENN1hGoEZAE/oTQvsVWK9lE1Sg1bnAXqeYknaSLXkxAnsk/qqdhsun
PINddjfPq0i7IaBvSkeT4/VpWhxADrQ9DHd2JUTBDpOzeIbjNYPNhdQoaUBjKn3z
n2B1CeKL+1DvZb4vxj0jKtAb78dYWqppVZ+TY6mMnxJFjIIKfhFclyLpzRPnhIN2
ibtX5qXNUHhVYgMsbXYkF8ejEbTWxza3LCKd5hHmCoHP6bmD+BHejMFl33e5YEHs
0snu2JndkpuU+BWH7ZM/lTmDpnjLPlmVZb4V106kaCmkwNdVwmIyOSFrs0eXhDJL
1f33emtLInit8832yCUMDG8nM0DVrX4niJWdpmS+ZWyeTdNRB/Bw+kpCWTOqEO/5
jp9y24x2DVfEF56cvZ/w2rJeG4NJg8a4nSI5t6/f0zaGatVxOzDPSYB6W7HRw06j
dAdIIcsGZFpibP6A2n/LAekvsCbEqTh+foTXkLi7PQWctIJBSH6SX5WAyhzh3nHZ
o8WsEDM5wiGv3Nxo876AsLxBOsob5BV1eZqqTzuDF002fdB5koqmPUK2PvEWaHLg
5Myx5cYJj2lLHsH4LpWjKIrcmXVtp5JEiOL0cIEw6wBMwSA6GQeGKnK7fs4CnLxv
qPYZDNXHapAB4JUCQ579w+agzruHH/+bScsdFeI4gNrkpfwbDjRQIxXcbOjz8Gkn
FRETMBq+imr3BbTKpfLK7BJrgfEUCnfxaviop85jmd3bTMsSCW0t43kDxzz+xTP3
UCEN+CntgZGv0p7qHVTu6hm7y/NYm2Dxns+JjrrKxtQIcSBnHgpZIzf1E3VJ9d1d
p9mCjOM3dtBApQCd7gkZfiN0q9NLJ9bxsgZdpQoWk+tXucLFRru/2Pk/NiPr7jCe
GLLR92QAVFTdCnMmr/IhLXWwjg1cpS7/71b4cdwIm5iCvbd8KD4kg1rveRV2B3ov
5kSrx1Opvon9GW9z6rLKDnskjQcIOH66yJa6LrmF/QiYcU9lE+loexKFKjMVNv32
ZtByb5bUSL84sj3sv1Y9GDmI8CNl9leF4q7dlO6QOKBbkTSBBlN0QMwYOmv1eq3V
MQmSMH7oozhHfd/wMU3ThLTP9t64viOIebMqIeWp8e+HajhORMsi2Ca/T8OF6sHQ
duxGXnPqMVo83kN8mqUOaMeT0APBfHbE96QpcSRe49gvgDHVWS1ROFzKonCIPyDr
LxdvrFC8XVMfgCpTWaG2bAbYAAqcKKb/IijsxZVZqvaeHxbif8+0LWrQXcF91RJE
NZuqMeYMwXw+CIEj8ay/ypQjKfgsyNLp3CmDD26s0ardgvVXfvF5ouLb6wlh8oJ9
8fo4ShEdVoSqZ+o9qCWzG/j1xpV2K7CN7liVH2SFzAqttn/75Uo1JJGFR7pMqBCz
drDOrc/y9p5MxEcZ+OKK6mqFVNRq3ykECD63wN0O9NY4E38Q3kXZoL3Q2zDBYriS
LBE1pLlu7MCBasH63Sw4ukT3UgwbEmGALZurwgSOyKpl3eQSNnyb+pHFVBuZrs/C
EADcEeqv9G56mwNSToWzp7mZicOE4/jK18cYxJzpGZw/hu2lRvjTLlBVyxB7oNTn
SFqrnw29RcneW5Qa2F9PFh8yf4lZXahNyig0JZrIeREy6PQaoZha1kP9rFLRnS7R
mNIfObs4zdm+34eQ9HSLOXZV6Oi4SVMIhwsuOfi+6XhM4oI3+awXtCL31MQRC++a
4Y4crAIFF3Uoxf/OjDwh/rvyFMrPfFN14NVKGXDWAtcUWAlM9TvmiT6nqzELgNZk
zTGw377fnGvTZeWB3NERnu9mHfRFCA1E1EhsJR/bLGoqtgwyOJZQMdxX2xXenP7G
84m4xsq6RozUmC/ySMsLBmC0OQVnnEmxf+OSbfI3zsbMj7LAQAkAvM4eTCfmGDEr
xosRz+HnDDxVin0/qfCUp6YsYyR5SvaS7JL/e/aoDRkUN+1uEdi2FgzijsuFPcAn
9R59AjBSOtvS95970CPe5udq8l/5fRYe/2nXLX3Hai0wU1zSK2vHb2RUDx8DAp/C
XJigP+iqtIHQCk68vwcE3Fd/Veu5SYASTq55E+dCosFPuS0HnOQcETrlIR+lvscq
YvmwZS+btNqiv9i4I26Jz0Olh3WiL07B6zGCNZeAzFI+lTCDSxkLWqdg3I1yzCIl
ug0QGVMnzLJbgCPJvgIG13032mGaq4T+uullFN8uu770l0fAgHHfMSpBVseX/1XJ
yVnbWjGeVTlwBPgs7noMHp2JpQEyFmB0m6/XeHQtRyTswSe8WDOpStANwMgpz10S
F4ARZQ8lBtZl01Ekqx60wxi+vh04BhFmEcVTzNh4bAD34UwnvyEknSdVXM57y7Z9
+YxY8ZHj6AklH8iiOhc4YDtKRjkUvFBmOnTHDqkWIhk/+c1yV9rpqx3VHGTYJfj9
npeW71zVeNqsVtZ6vtaOU0gNqYY8z7LOdbjZ7eDbmVX+x6GfFz9+XRK2sA9UssF0
aKnatt5LPmqsDEUnOkRP+5WY4zPy/NecL929WmpOCODyy7pgxhMMD1c+ps2X/xTG
1Rd8SK3NEe3jvhftAIB4iYtlGQFEBylmP6PP3RqEEuQQzNFJGAhk3o8eCh/kfH7z
caoWHTtYtqNHfA391p7IC5Y7kq+NpKhUWW1Ab1hZLQ1F/LZUtTpMazp4ZLDehcoO
8te5ca+/4KCcaCyWOPflMUiMQ0HL2gd/DxL7VNcQSZlWLpUd/8e4JTA9q6JUSQGx
GUUGYnwHp/l3/m55XspCPhtCIVP8wIZMzivnYLnMtNm4s3RYU93RMPVuidkQD5Uf
8gj8lvvpQqbrxfAXV1HGhks2BIqodi/fpE++2mRQ7EhZgCbP+PxoImdIFzHxgY7X
WPDN5D4edJB0kk9gaBeWLicNiiu3PUiK4NTJnEI0QPjRjmbU0mEEhuGpKR94hQCr
mM2W8CGccn4MQ0/Gwg6sgIcU10CETXbAIVXIMqiXJU/ICG+BOBxFSkN3LqR3BflJ
Z+HjlE+0E1GHVJkqB0iRLup6LOuON6ddzc0k3o0PEcpqoUkNDmyW/s+CtvQGP2PD
f20+HfgxoUI5BnyXpxvdCoUfAgSA7Ev1sMrJHorOuIaBSOoDIujszLr0x39m+UAn
tF9K3cPhXJJvbwUGC75sGMivAsEDE13ZkqQNTvxcA6WD7wc8tLD5DzZG2gqjNPGu
vZ9WPErxXn0UtZ89wx8rO0i+TJ5AT+uGRfkcDmSPnklG1AmgL1fccV0d6dyk0hkV
PrGfUlCFOwcZUKDAE1ZSez9chX9EcKUZcwIunJuy8jRKnXMt9O+lvUHF65zZXIxS
HlCTzqImIeWitYxmRn8h9C8LyZt3w2WzXb3CCAdJFJqV87HaBQibSQKoDFTYsJ4Y
LYOlmHS3gl+BFtbXXoC+OmVewW0NVYmTcjnIP2oGsLqHmqZjqFmR2hvPd5/zEPns
NspMshIsYZA+XtOfKpn/Uqph9Ceg4rTNlMLtrnlwI7d5XgaHDwxFqsX3+f+vfuyt
KAOtojI7ygX2CxpGycqLssmwSJkv0RC8IHoeQ8HLrWFjGqC/DnTsXBjuAxJFiXmN
QSymc74b+J7UKqTHGhtt/cXJXlsm0kvA9Q1npPSCe+qZDdPKf9YiT+zj4HUoRF4X
wIKb5iACuKI7zlO0vi9kISQVz7NJFvMEWz14FBYCcPsyNMIMu4la3g2IE37+gj95
NvkAPaagBdF20NMnjXlnFXAXAPfpoDGfAWtV7qurlstQZp5PSvsjL6ef6q0dKZz2
HehKYbxJZ3fXo5xeOeD2iKuEsldg9tJesY67kbHkwrX0VvxxmooOdjpg1IOFDLaf
ikQn9fe+PKlgk054nU+C94++IusKABR/ZUHw3ZqNR0pC/OtDqBQCKeIIUeZU6CH2
b7Fj+HyfSnc5hn2RFLzB8VSQM/ox+8E5uRZMHdDfH+FsKP6T2UC4tnQJALf29uan
pH8td/M4m/YZ7os3I4jdYJPPi+76sRvHwYLLnWKw+AOyZQKhgTlHvVhac68bVtIi
fWOCilJeaS34vhrQhe7mgQROeqG2lHawR4sdUqdGGZPQgVhYdMcGCKlS8dtS7csp
d1yKtLqg/vp+XbuUppr9Rp/segZW/9aaXcqrplSx9uNiIPXSqNi8+8MtTejYjB7t
A1PVeAiiL9w6zBS2mKwGJf31DrIyKS0zwD9K7CwZZDwDQuAEpnHlS5SAgCF3lPcY
SmHNkaoY/RZ05ZcJ5YxHoGHv8RGZ6aTzjvS6bQ52dMMr9tzdQH9qATb+4uou4Rk5
2baNUf2MHVE1O0Cds/m5uTVzI5uW9LsJC1yLXC3LAvXBsXHRDPgZ+1kemKBlExOj
cNw9uw5OCV/zxaMpEE3fIAWVSWaZqiOuae3KWpYdmA3yF6krHpyGrnLk9YaEIypl
8s9ExxS0NeanFrskfi105C8FrttW2iPRxGHinpctuD/EFHnhVFW3c+QmlsNAYjAk
mJZCwwdyBfxqBn9/CgPhRKdiuOU8kkDf1+gGydngprwrTbBYJWFt12mInLXr3e/B
gw0X5nRPAaRue5oGMgHj6VsrL46k7bUQ8gijsXpwNuuiklwttXMeYPM5h+UJkY2B
jQClnjvfC1E2+OEEYyDJhbYWVRV2ei8LTxrFNYZTBbiYWE4dScgODcGyHQS6Mm7A
tALS/CNv59knV76d0TlrjFmvwbgJeL9bLbdReo11ZHe/XZrsYu8XpwvcG95mjiqO
2eRXCF4lUH/pZCLMPuyp+ElN8eLkv3jLBwFEXEHAElAtrcDPuZPuAWP1FOL+aDlI
O1PpE784BE35Hh+Km6r7yxEhi/LxfttVi1jVb5iek6kj+07QMG0nI/T9LReR03ew
zTWl3lyzMv97GWlL3VOMH8TbhQTsaw0S/Y/KqyaQxvGViRuGNoZylcxScd4G83hc
xPGfBQgFeMKaj7/Pb6mJ8MKDu1Pwe8lUQP8h2MIvF8FmqOD0T/qLUkaMvv21l/j3
1FI46FGOtUOwkhka+jNJtoWJKgXwr3h9fn46iWfhk+7+g+RBJLIGl6inPzW0R0v4
GpLnDDBqiyW9bSAIIUpn076DCUC5Y1LCmDZe8hb/iR1rksfDoZFHEw+MYRqMZMh+
5kOLLkPQ6yRYKABfCsYOE8Vq8YsSDN+g+JI5qED71Ly4AIq+VS4/L0H6DG3KUcSq
9oFAD91z1E159Kj6C1XxLRcYOU9QxGCyNXwdnkAQwb/pquE2zuqwqjCO6PzdRzRh
RD6xEPeitnDF3o7U2w5p3rDjnzzPGXVBnm5hg9oi8AYvHqIlQKIqH2QcDFOgMudY
IXAspxLiRhjZ3SGqtMyJvIUAqR5VAllwSiGhaK9J00kT0TiaHsylOspWxWmYwye7
r+JP1UcSrbaQcS6PbtOmVQ8embfq74mjvaSjrIhKa7S5mBGW3IcXoSDLjboDZTtq
7zwF7nUPEEZ25S2yHyZqke0yDHiWM80Q3WcDYnIYL2xuE1LGgpMtMhfz8J5svudG
32eX2Tl0ZVqsjPU06GsVEz2EF9UgPM9zpjAWPIW9e0GEP7crY82hg1Ji7GtD0acP
KWAu34jaOrgtUtx1mX0xTbNszqkD1Md3IZHipDcVPyS65q6ztO9hsI1gTvwFehLR
ozbT+R5cAFTmRval7+V7OhIhkfo7M61PTOELvElXJHZ+G6ehOSw/jJsSPRoMl760
WAv4dWhIAY3xpcpV77zwR8Nw8UPFOo/VGfypqtMtNIE2I+SCxYns88Oq6VEsAWmK
RbHPu4ngiLZyfrP+AsDa831f2Ct70yeAetN0Y3gBMxRcLCbqO6V2oYpEmMC9zBgX
h5AUzQKNruGDBZg3l39nfKOtXibjoIYZMR2QxRiczTgsaX0tfdk7JD3F7Xdt1Z7i
oZGTS+wksOvSMXGNGkwd+x5QZNvAk/M2OAntkAB8/Ry/z48KSwRxPjNyUsHkr4VG
gywBHfTIEx3dKLkd6ADcbyuFZMWqE4s4IBSJclrC8r6PNIXAYSfzzMMswAYHw7BS
tlj8GBFWdRL4pJaQKIZA2rH+hWGlE+e44WokL9zgVCKtoeWeLPyGz5fFABZoK6uf
BTB8ZBtQfTlFWmMQ7/4+bRgQm2qT+6owBkeWQ78B7OwXHLYrhL3ZKeKxsVbkqJJb
f3VHhhfIThpU5ALbE7HDvRoJo7Qxib4w5g4wb93wMxN4Jm0iiTlQmmFZ2cvhRmak
bwCYcnKGYw0Fxp8E1KCsB/kfcrMjKhfDaWTQkwG9hJxGcozEt5PQnq0S2dnfsU5b
vqAg7GTG6bZdNyaTcHevMVkiOQ3fKrJJ0/7zI0zlNA5jMcnGfU7TVxtkiwWJmY1s
6i7hjUoMC4Wk3MRdvU/QRkxfz+SO/zYorWdUb4cKvYxx3QsdWn2TQSULt2jwgMoh
hE9XaII9DpY/Ao2Mc+5k45oUmmQluhBbXkhHKh1i2ESB4xi/LiyGGXpqDz969L8C
XGu26i0gE3Z7D6Gnf1FUQ92S9tmw5Uzed8+R2Nt+01RgtbHR/sUjcnZe/gjYi0JW
OlxKdFxK+v2vFpRmlnCxadmunS1f/su+C15GE2Irl8AOAgO8eUdCyngpT4Y3uueD
v1rjXdKPd5fHq/Sq+oQ5gM5GFf+Ne0KtN2KH3+9Nw7hsZS/7Dhi78RoB8K0+4PNv
nMfW5FRATP7eHSzDZP0vuE90yinL3NjMEkB7P5/dEp1OwHI7GEx/6k10zex0DpM5
SMjPHM+PLAKHovQpZPHzyE8zmqS1FmXANSPy7ShhYmSGczWex+zMJtiOkvdVCklT
jl9uIx5C6mg8xRJy6gt7YdKvnsUfiD5Z/h9wA4jmlDLV1kTbZWlS8tU3Y2+wqrZ+
5ZJSXw84rl70eleWs10B9jqyQhQKDOLqHupYARcQViM=
`pragma protect end_protected

//pragma protect end
