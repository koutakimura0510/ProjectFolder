/*
 * Create 2022/4/21
 * Author koutakimura
 * -
 * 独自バスシステムのラッパーモジュール
 */
module usibWrapper (
    input           iClk,      // バスシステムのクロック指定
    input           iRst       // Active High
);



endmodule