/*-----------------------------------------------------------------------------
 * Create  2023/4/13
 * Author  koutakimura
 * -
 * シンセサイザーの制御を行う。
 * MIDI 信号をデコードし、パラメータ設定に則ってサウンドを生成する。
 * 
 * V1.0 new release
 *-----------------------------------------------------------------------------*/
module SynthesizerUnit (
	// AUDIO OUT
	output [31:0] oAUDIO,
    // CLK Reset
	input  iMRST,
    input  iSRST,
	input  iMCLK,
    input  iSCLK
);





endmodule