//----------------------------------------------------------
// Create 2022/4/21
// Author koutakimura
// -
// 独自バスシステムのラッパーモジュール
// 
// ID | module
// ----------------------
// 01 | PFBWrapper
// 02 | ~~~~
// 03 | ~~~~
// 
// 上記のようにモジュールを ID で振り分ける
// 各モジュールに CSR (コントロール・ステータスレジスタ) を作成し、
// Bus を経由して、
// if (!ID) などと、IDが異なっていたらスルーするようにする。
// 
//----------------------------------------------------------
module usibWrapper (
    input           iClk,      // バスシステムのクロック指定
    input           iRst       // Active High
);



endmodule