
//
// Verific Verilog Description of module MTopTi180MIPI25GRxHDMIV101
//

module MTopTi180MIPI25GRxHDMIV101 (MipiDphyRx1_RESET_N, MipiDphyRx1_RST0_N, 
            MipiDphyRx1_STOPSTATE_CLK, MipiDphyRx1_STOPSTATE_LAN0, MipiDphyRx1_STOPSTATE_LAN1, 
            MipiDphyRx1_ERR_ESC_LAN0, MipiDphyRx1_ERR_ESC_LAN1, MipiDphyRx1_ERR_CONTROL_LAN0, 
            MipiDphyRx1_ERR_CONTROL_LAN1, MipiDphyRx1_TX_REQUEST_ESC, MipiDphyRx1_TURN_REQUEST, 
            MipiDphyRx1_FORCE_RX_MODE, MipiDphyRx1_TX_TRIGGER_ESC, MipiDphyRx1_RX_TRIGGER_ESC, 
            MipiDphyRx1_DIRECTION, MipiDphyRx1_ERR_CONTENTION_LP0, MipiDphyRx1_ERR_CONTENTION_LP1, 
            MipiDphyRx1_RX_CLK_ACTIVE_HS, MipiDphyRx1_RX_ACTIVE_HS_LAN0, 
            MipiDphyRx1_RX_ACTIVE_HS_LAN1, MipiDphyRx1_RX_VALID_HS_LAN0, 
            MipiDphyRx1_RX_VALID_HS_LAN1, MipiDphyRx1_RX_SYNC_HS_LAN0, MipiDphyRx1_RX_SYNC_HS_LAN1, 
            MipiDphyRx1_RX_SKEW_CAL_HS_LAN0, MipiDphyRx1_RX_SKEW_CAL_HS_LAN1, 
            MipiDphyRx1_RX_DATA_HS_LAN0, MipiDphyRx1_RX_DATA_HS_LAN1, MipiDphyRx1_ERR_SOT_HS_LAN0, 
            MipiDphyRx1_ERR_SOT_HS_LAN1, MipiDphyRx1_ERR_SOT_SYNC_HS_LAN0, 
            MipiDphyRx1_ERR_SOT_SYNC_HS_LAN1, MipiDphyRx1_RX_LPDT_ESC, MipiDphyRx1_RX_DATA_ESC, 
            MipiDphyRx1_RX_VALID_ESC, MipiDphyRx1_RX_ERR_SYNC_ESC, MipiDphyRx1_TX_LPDT_ESC, 
            MipiDphyRx1_TX_DATA_ESC, MipiDphyRx1_TX_VALID_ESC, MipiDphyRx1_TX_READY_ESC, 
            MipiDphyRx1_TX_ULPS_ESC, MipiDphyRx1_TX_ULPS_EXIT, MipiDphyRx1_RX_ULPS_CLK_NOT, 
            MipiDphyRx1_RX_ULPS_ACTIVE_CLK_NOT, MipiDphyRx1_RX_ULPS_ESC_LAN0, 
            MipiDphyRx1_RX_ULPS_ESC_LAN1, MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN0, 
            MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN1, MipiDphyRx1_WORD_CLKOUT_HS, 
            MipiDphyRx1_LP_CLK, MipiDphyRx1_RX_CLK_ESC_LAN0, MipiDphyRx1_RX_CLK_ESC_LAN1, 
            MipiDphyRx1_TX_CLK_ESC, oAdv7511Vs, oAdv7511Hs, oAdv7511De, 
            oAdv7511Data, iAdv7511Sda, oAdv7511SdaOe, iAdv7511Scl, oAdv7511SclOe, 
            oLed, iPushSw, iSCLK, iBCLK, iPCLK, iFCLK, pll_inst1_LOCKED, 
            pll_inst1_RSTN, iVCLK, pll_inst2_LOCKED, pll_inst2_RSTN, 
            oTestPort, jtag_inst1_TDI, jtag_inst1_TCK, jtag_inst1_TMS, 
            jtag_inst1_TDO, jtag_inst1_SEL, jtag_inst1_DRCK, jtag_inst1_RUNTEST, 
            jtag_inst1_CAPTURE, jtag_inst1_SHIFT, jtag_inst1_UPDATE, jtag_inst1_RESET, 
            jtag_inst2_CAPTURE, jtag_inst2_DRCK, jtag_inst2_RESET, jtag_inst2_RUNTEST, 
            jtag_inst2_SEL, jtag_inst2_SHIFT, jtag_inst2_TCK, jtag_inst2_TDI, 
            jtag_inst2_TMS, jtag_inst2_UPDATE, jtag_inst2_TDO);
    output MipiDphyRx1_RESET_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_RST0_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_STOPSTATE_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTROL_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTROL_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_REQUEST_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TURN_REQUEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_FORCE_RX_MODE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [3:0]MipiDphyRx1_TX_TRIGGER_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [3:0]MipiDphyRx1_RX_TRIGGER_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_DIRECTION /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTENTION_LP0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_CONTENTION_LP1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ACTIVE_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ACTIVE_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ACTIVE_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SYNC_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SKEW_CAL_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_SKEW_CAL_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_ERR_SOT_SYNC_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_LPDT_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]MipiDphyRx1_RX_DATA_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_VALID_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ERR_SYNC_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_LPDT_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]MipiDphyRx1_TX_DATA_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_VALID_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_READY_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_ULPS_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output MipiDphyRx1_TX_ULPS_EXIT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_CLK_NOT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_CLK_NOT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_ULPS_ACTIVE_NOT_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_WORD_CLKOUT_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_LP_CLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input MipiDphyRx1_RX_CLK_ESC_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output MipiDphyRx1_TX_CLK_ESC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511Vs /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511Hs /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output oAdv7511De /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [15:0]oAdv7511Data /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iAdv7511Sda /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output oAdv7511SdaOe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iAdv7511Scl /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output oAdv7511SclOe /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [5:0]oLed /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [1:0]iPushSw /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iSCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iBCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iPCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input iFCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_inst1_LOCKED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output pll_inst1_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input iVCLK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_inst2_LOCKED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output pll_inst2_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [25:0]oTestPort /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst2_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst2_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    
    wire la0_probe10, la0_probe2, rFRST, rBRST, rVRST, rnVRST, la0_probe11, 
        \la0_probe6[0] , \la0_probe9[0] , \MCsiRxController/MCsi2Decoder/rHsSt[0] , 
        \la0_probe3[0] , \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd , 
        la0_probe4, la0_probe5, la0_probe7, n116, n117, la0_probe0, 
        n119, n120, \MCsiRxController/wHsPixel[0] , \MCsiRxController/MCsi2Decoder/wFtiRvd[0] , 
        wCddFifoFull, n124, n125, \MCsiRxController/wHsValid , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] , 
        \MCsiRxController/MCsi2Decoder/rHsSt[2] , \MCsiRxController/MCsi2Decoder/rHsSt[1] , 
        \la0_probe9[7] , \la0_probe9[6] , \la0_probe9[5] , \la0_probe9[4] , 
        \la0_probe9[3] , \la0_probe9[2] , \la0_probe9[1] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] , 
        \MCsiRxController/MCsi2Decoder/wFtiEmp[0] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
        n169, n170, \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[16] , n189, n190, \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9] , 
        n210, n211, \MCsiRxController/wHsPixel[1] , \MCsiRxController/wHsPixel[2] , 
        \MCsiRxController/wHsPixel[3] , \MCsiRxController/wHsPixel[4] , 
        \MCsiRxController/wHsPixel[5] , \MCsiRxController/wHsPixel[6] , 
        \MCsiRxController/wHsPixel[7] , \MCsiRxController/wHsPixel[8] , 
        \MCsiRxController/wHsPixel[9] , \MCsiRxController/wHsPixel[10] , 
        \MCsiRxController/wHsPixel[11] , \MCsiRxController/wHsPixel[12] , 
        \MCsiRxController/wHsPixel[13] , \MCsiRxController/wHsPixel[14] , 
        \MCsiRxController/wHsPixel[15] , \wHsWordCnt[1] , \wHsWordCnt[2] , 
        \wHsWordCnt[3] , \wHsWordCnt[4] , \wHsWordCnt[5] , \wHsWordCnt[6] , 
        \wHsWordCnt[7] , \wHsWordCnt[8] , \wHsWordCnt[9] , \wHsWordCnt[10] , 
        \wHsWordCnt[11] , \wHsWordCnt[12] , \wHsWordCnt[13] , \wHsWordCnt[14] , 
        \wHsWordCnt[15] , \wHsDatatype[2] , \wHsDatatype[3] , \wHsDatatype[4] , 
        \wHsDatatype[5] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] , \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] , 
        \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] , \la0_probe8[0] , 
        \la0_probe8[1] , \la0_probe8[2] , \la0_probe8[3] , \la0_probe8[4] , 
        \la0_probe8[5] , \la0_probe8[6] , \la0_probe8[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] , wVideoVd, n295, 
        n296, \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] , \MCsiRxController/wFtiEmp[0] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] , 
        \wVideoPixel[0] , \wVideoPixel[1] , \wVideoPixel[2] , \wVideoPixel[3] , 
        \wVideoPixel[4] , \wVideoPixel[5] , \wVideoPixel[6] , \wVideoPixel[7] , 
        \wVideoPixel[8] , \wVideoPixel[9] , \wVideoPixel[10] , \wVideoPixel[11] , 
        \wVideoPixel[12] , \wVideoPixel[13] , \wVideoPixel[14] , \wVideoPixel[15] , 
        n331, n332, \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] , 
        \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] , 
        \la0_probe6[1] , \la0_probe6[2] , \la0_probe6[3] , \la0_probe6[4] , 
        \la0_probe6[5] , \la0_probe6[6] , \la0_probe6[7] , \la0_probe6[8] , 
        \la0_probe6[9] , \la0_probe6[10] , \la0_probe6[11] , \la0_probe6[12] , 
        \la0_probe6[13] , \la0_probe6[14] , \la0_probe6[15] , \la0_probe3[1] , 
        \MVideoPostProcess/rVtgRstCnt[0] , \MVideoPostProcess/rVtgRST[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] , \MVideoPostProcess/inst_adv7511_config/r_m_en_1P , 
        \MVideoPostProcess/inst_adv7511_config/r_last_1P , \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] , \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P , \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] , 
        \MVideoPostProcess/inst_adv7511_config/w_ack , \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] , n436, n437, 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] , 
        \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] , \MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] , 
        \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] , \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] , \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] , 
        \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] , 
        \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] , \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] , 
        \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] , 
        n489, n490, \MVideoPostProcess/mVideoTimingGen/rVpos[0] , n492, 
        n493, \MVideoPostProcess/mVideoTimingGen/rVde[0] , \MVideoPostProcess/mVideoTimingGen/rHpos[0] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[1] , \MVideoPostProcess/mVideoTimingGen/rVpos[2] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[3] , \MVideoPostProcess/mVideoTimingGen/rVpos[4] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[5] , \MVideoPostProcess/mVideoTimingGen/rVpos[6] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[7] , \MVideoPostProcess/mVideoTimingGen/rVpos[8] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[9] , \MVideoPostProcess/mVideoTimingGen/rVpos[10] , 
        \MVideoPostProcess/mVideoTimingGen/rVpos[11] , \MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre , 
        \MVideoPostProcess/mVideoTimingGen/rVde[1] , \MVideoPostProcess/mVideoTimingGen/rVde[3] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[1] , \MVideoPostProcess/mVideoTimingGen/rHpos[2] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[3] , \MVideoPostProcess/mVideoTimingGen/rHpos[4] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[5] , \MVideoPostProcess/mVideoTimingGen/rHpos[6] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[7] , \MVideoPostProcess/mVideoTimingGen/rHpos[8] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[9] , \MVideoPostProcess/mVideoTimingGen/rHpos[10] , 
        \MVideoPostProcess/mVideoTimingGen/rHpos[11] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] , 
        wVideofull, n532, n533, \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] , 
        n555, n556, \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] , 
        n573, n574, \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] , 
        n596, n597, \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] , 
        n614, n615, \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] , 
        n637, n638, \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] , 
        n655, n656, \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] , 
        n678, \MVideoPostProcess/rVtgRstCnt[1] , \MVideoPostProcess/rVtgRstCnt[2] , 
        \MVideoPostProcess/rVtgRstCnt[3] , \MVideoPostProcess/rVtgRstCnt[4] , 
        \MVideoPostProcess/rVtgRstCnt[5] , \MVideoPostProcess/rVtgRstCnt[6] , 
        \MVideoPostProcess/rVtgRstCnt[7] , \MVideoPostProcess/rVtgRstCnt[8] , 
        \MVideoPostProcess/rVtgRstCnt[9] , \MVideoPostProcess/rVtgRstCnt[10] , 
        \MVideoPostProcess/rVtgRST[1] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] , 
        \genblk1.genblk1[0].mPulseGenerator/rSft[0] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] , 
        \genblk1.genblk1[0].mPulseGenerator/rSft[1] , \genblk1.genblk1[0].mPulseGenerator/rSft[2] , 
        \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] , \genblk1.genblk1[1].mPulseGenerator/rSft[0] , 
        \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] , \genblk1.genblk1[1].mPulseGenerator/rSft[1] , 
        \genblk1.genblk1[1].mPulseGenerator/rSft[2] , \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] , 
        \genblk1.genblk1[3].mPulseGenerator/rSft[0] , \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] , 
        \genblk1.genblk1[3].mPulseGenerator/rSft[1] , \genblk1.genblk1[3].mPulseGenerator/rSft[2] , 
        \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] , \genblk1.genblk1[4].mPulseGenerator/rSft[0] , 
        \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] , \genblk1.genblk1[4].mPulseGenerator/rSft[1] , 
        \genblk1.genblk1[4].mPulseGenerator/rSft[2] , \edb_top_inst/n2759 , 
        \edb_top_inst/la0/la_run_trig , \edb_top_inst/la0/la_trig_pattern[0] , 
        \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig , 
        \edb_top_inst/la0/la_capture_pattern[0] , \edb_top_inst/la0/la_trig_mask[0] , 
        \edb_top_inst/la0/la_num_trigger[0] , \edb_top_inst/la0/la_window_depth[0] , 
        \edb_top_inst/la0/la_soft_reset_in , \edb_top_inst/la0/address_counter[0] , 
        \edb_top_inst/la0/opcode[0] , \edb_top_inst/la0/bit_count[0] , \edb_top_inst/la0/word_count[0] , 
        \edb_top_inst/la0/data_out_shift_reg[0] , \edb_top_inst/la0/module_state[0] , 
        \edb_top_inst/la0/la_resetn_p1 , \edb_top_inst/la0/la_resetn , \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/cap_fifo_din_cu[0] , \edb_top_inst/la0/cap_fifo_din_tu[0] , 
        \edb_top_inst/la0/internal_register_select[0] , \edb_top_inst/la0/la_trig_pos[0] , 
        \edb_top_inst/la0/la_trig_pattern[1] , \edb_top_inst/la0/la_capture_pattern[1] , 
        \edb_top_inst/la0/la_trig_mask[1] , \edb_top_inst/la0/la_trig_mask[2] , 
        \edb_top_inst/la0/la_trig_mask[3] , \edb_top_inst/la0/la_trig_mask[4] , 
        \edb_top_inst/la0/la_trig_mask[5] , \edb_top_inst/la0/la_trig_mask[6] , 
        \edb_top_inst/la0/la_trig_mask[7] , \edb_top_inst/la0/la_trig_mask[8] , 
        \edb_top_inst/la0/la_trig_mask[9] , \edb_top_inst/la0/la_trig_mask[10] , 
        \edb_top_inst/la0/la_trig_mask[11] , \edb_top_inst/la0/la_trig_mask[12] , 
        \edb_top_inst/la0/la_trig_mask[13] , \edb_top_inst/la0/la_trig_mask[14] , 
        \edb_top_inst/la0/la_trig_mask[15] , \edb_top_inst/la0/la_trig_mask[16] , 
        \edb_top_inst/la0/la_trig_mask[17] , \edb_top_inst/la0/la_trig_mask[18] , 
        \edb_top_inst/la0/la_trig_mask[19] , \edb_top_inst/la0/la_trig_mask[20] , 
        \edb_top_inst/la0/la_trig_mask[21] , \edb_top_inst/la0/la_trig_mask[22] , 
        \edb_top_inst/la0/la_trig_mask[23] , \edb_top_inst/la0/la_trig_mask[24] , 
        \edb_top_inst/la0/la_trig_mask[25] , \edb_top_inst/la0/la_trig_mask[26] , 
        \edb_top_inst/la0/la_trig_mask[27] , \edb_top_inst/la0/la_trig_mask[28] , 
        \edb_top_inst/la0/la_trig_mask[29] , \edb_top_inst/la0/la_trig_mask[30] , 
        \edb_top_inst/la0/la_trig_mask[31] , \edb_top_inst/la0/la_trig_mask[32] , 
        \edb_top_inst/la0/la_trig_mask[33] , \edb_top_inst/la0/la_trig_mask[34] , 
        \edb_top_inst/la0/la_trig_mask[35] , \edb_top_inst/la0/la_trig_mask[36] , 
        \edb_top_inst/la0/la_trig_mask[37] , \edb_top_inst/la0/la_trig_mask[38] , 
        \edb_top_inst/la0/la_trig_mask[39] , \edb_top_inst/la0/la_trig_mask[40] , 
        \edb_top_inst/la0/la_trig_mask[41] , \edb_top_inst/la0/la_trig_mask[42] , 
        \edb_top_inst/la0/la_trig_mask[43] , \edb_top_inst/la0/la_trig_mask[44] , 
        \edb_top_inst/la0/la_trig_mask[45] , \edb_top_inst/la0/la_trig_mask[46] , 
        \edb_top_inst/la0/la_trig_mask[47] , \edb_top_inst/la0/la_trig_mask[48] , 
        \edb_top_inst/la0/la_trig_mask[49] , \edb_top_inst/la0/la_trig_mask[50] , 
        \edb_top_inst/la0/la_trig_mask[51] , \edb_top_inst/la0/la_trig_mask[52] , 
        \edb_top_inst/la0/la_trig_mask[53] , \edb_top_inst/la0/la_trig_mask[54] , 
        \edb_top_inst/la0/la_trig_mask[55] , \edb_top_inst/la0/la_trig_mask[56] , 
        \edb_top_inst/la0/la_trig_mask[57] , \edb_top_inst/la0/la_trig_mask[58] , 
        \edb_top_inst/la0/la_trig_mask[59] , \edb_top_inst/la0/la_trig_mask[60] , 
        \edb_top_inst/la0/la_trig_mask[61] , \edb_top_inst/la0/la_trig_mask[62] , 
        \edb_top_inst/la0/la_trig_mask[63] , \edb_top_inst/la0/la_num_trigger[1] , 
        \edb_top_inst/la0/la_num_trigger[2] , \edb_top_inst/la0/la_num_trigger[3] , 
        \edb_top_inst/la0/la_num_trigger[4] , \edb_top_inst/la0/la_num_trigger[5] , 
        \edb_top_inst/la0/la_num_trigger[6] , \edb_top_inst/la0/la_num_trigger[7] , 
        \edb_top_inst/la0/la_num_trigger[8] , \edb_top_inst/la0/la_num_trigger[9] , 
        \edb_top_inst/la0/la_num_trigger[10] , \edb_top_inst/la0/la_num_trigger[11] , 
        \edb_top_inst/la0/la_num_trigger[12] , \edb_top_inst/la0/la_num_trigger[13] , 
        \edb_top_inst/la0/la_num_trigger[14] , \edb_top_inst/la0/la_num_trigger[15] , 
        \edb_top_inst/la0/la_num_trigger[16] , \edb_top_inst/la0/la_window_depth[1] , 
        \edb_top_inst/la0/la_window_depth[2] , \edb_top_inst/la0/la_window_depth[3] , 
        \edb_top_inst/la0/la_window_depth[4] , \edb_top_inst/la0/address_counter[1] , 
        \edb_top_inst/la0/address_counter[2] , \edb_top_inst/la0/address_counter[3] , 
        \edb_top_inst/la0/address_counter[4] , \edb_top_inst/la0/address_counter[5] , 
        \edb_top_inst/la0/address_counter[6] , \edb_top_inst/la0/address_counter[7] , 
        \edb_top_inst/la0/address_counter[8] , \edb_top_inst/la0/address_counter[9] , 
        \edb_top_inst/la0/address_counter[10] , \edb_top_inst/la0/address_counter[11] , 
        \edb_top_inst/la0/address_counter[12] , \edb_top_inst/la0/address_counter[13] , 
        \edb_top_inst/la0/address_counter[14] , \edb_top_inst/la0/address_counter[15] , 
        \edb_top_inst/la0/address_counter[16] , \edb_top_inst/la0/address_counter[17] , 
        \edb_top_inst/la0/address_counter[18] , \edb_top_inst/la0/address_counter[19] , 
        \edb_top_inst/la0/address_counter[20] , \edb_top_inst/la0/address_counter[21] , 
        \edb_top_inst/la0/address_counter[22] , \edb_top_inst/la0/address_counter[23] , 
        \edb_top_inst/la0/address_counter[24] , \edb_top_inst/la0/address_counter[25] , 
        \edb_top_inst/la0/address_counter[26] , \edb_top_inst/la0/opcode[1] , 
        \edb_top_inst/la0/opcode[2] , \edb_top_inst/la0/opcode[3] , \edb_top_inst/la0/bit_count[1] , 
        \edb_top_inst/la0/bit_count[2] , \edb_top_inst/la0/bit_count[3] , 
        \edb_top_inst/la0/bit_count[4] , \edb_top_inst/la0/bit_count[5] , 
        \edb_top_inst/la0/word_count[1] , \edb_top_inst/la0/word_count[2] , 
        \edb_top_inst/la0/word_count[3] , \edb_top_inst/la0/word_count[4] , 
        \edb_top_inst/la0/word_count[5] , \edb_top_inst/la0/word_count[6] , 
        \edb_top_inst/la0/word_count[7] , \edb_top_inst/la0/word_count[8] , 
        \edb_top_inst/la0/word_count[9] , \edb_top_inst/la0/word_count[10] , 
        \edb_top_inst/la0/word_count[11] , \edb_top_inst/la0/word_count[12] , 
        \edb_top_inst/la0/word_count[13] , \edb_top_inst/la0/word_count[14] , 
        \edb_top_inst/la0/word_count[15] , \edb_top_inst/la0/data_out_shift_reg[1] , 
        \edb_top_inst/la0/data_out_shift_reg[2] , \edb_top_inst/la0/data_out_shift_reg[3] , 
        \edb_top_inst/la0/data_out_shift_reg[4] , \edb_top_inst/la0/data_out_shift_reg[5] , 
        \edb_top_inst/la0/data_out_shift_reg[6] , \edb_top_inst/la0/data_out_shift_reg[7] , 
        \edb_top_inst/la0/data_out_shift_reg[8] , \edb_top_inst/la0/data_out_shift_reg[9] , 
        \edb_top_inst/la0/data_out_shift_reg[10] , \edb_top_inst/la0/data_out_shift_reg[11] , 
        \edb_top_inst/la0/data_out_shift_reg[12] , \edb_top_inst/la0/data_out_shift_reg[13] , 
        \edb_top_inst/la0/data_out_shift_reg[14] , \edb_top_inst/la0/data_out_shift_reg[15] , 
        \edb_top_inst/la0/data_out_shift_reg[16] , \edb_top_inst/la0/data_out_shift_reg[17] , 
        \edb_top_inst/la0/data_out_shift_reg[18] , \edb_top_inst/la0/data_out_shift_reg[19] , 
        \edb_top_inst/la0/data_out_shift_reg[20] , \edb_top_inst/la0/data_out_shift_reg[21] , 
        \edb_top_inst/la0/data_out_shift_reg[22] , \edb_top_inst/la0/data_out_shift_reg[23] , 
        \edb_top_inst/la0/data_out_shift_reg[24] , \edb_top_inst/la0/data_out_shift_reg[25] , 
        \edb_top_inst/la0/data_out_shift_reg[26] , \edb_top_inst/la0/data_out_shift_reg[27] , 
        \edb_top_inst/la0/data_out_shift_reg[28] , \edb_top_inst/la0/data_out_shift_reg[29] , 
        \edb_top_inst/la0/data_out_shift_reg[30] , \edb_top_inst/la0/data_out_shift_reg[31] , 
        \edb_top_inst/la0/data_out_shift_reg[32] , \edb_top_inst/la0/data_out_shift_reg[33] , 
        \edb_top_inst/la0/data_out_shift_reg[34] , \edb_top_inst/la0/data_out_shift_reg[35] , 
        \edb_top_inst/la0/data_out_shift_reg[36] , \edb_top_inst/la0/data_out_shift_reg[37] , 
        \edb_top_inst/la0/data_out_shift_reg[38] , \edb_top_inst/la0/data_out_shift_reg[39] , 
        \edb_top_inst/la0/data_out_shift_reg[40] , \edb_top_inst/la0/data_out_shift_reg[41] , 
        \edb_top_inst/la0/data_out_shift_reg[42] , \edb_top_inst/la0/data_out_shift_reg[43] , 
        \edb_top_inst/la0/data_out_shift_reg[44] , \edb_top_inst/la0/data_out_shift_reg[45] , 
        \edb_top_inst/la0/data_out_shift_reg[46] , \edb_top_inst/la0/data_out_shift_reg[47] , 
        \edb_top_inst/la0/data_out_shift_reg[48] , \edb_top_inst/la0/data_out_shift_reg[49] , 
        \edb_top_inst/la0/data_out_shift_reg[50] , \edb_top_inst/la0/data_out_shift_reg[51] , 
        \edb_top_inst/la0/data_out_shift_reg[52] , \edb_top_inst/la0/data_out_shift_reg[53] , 
        \edb_top_inst/la0/data_out_shift_reg[54] , \edb_top_inst/la0/data_out_shift_reg[55] , 
        \edb_top_inst/la0/data_out_shift_reg[56] , \edb_top_inst/la0/data_out_shift_reg[57] , 
        \edb_top_inst/la0/data_out_shift_reg[58] , \edb_top_inst/la0/data_out_shift_reg[59] , 
        \edb_top_inst/la0/data_out_shift_reg[60] , \edb_top_inst/la0/data_out_shift_reg[61] , 
        \edb_top_inst/la0/data_out_shift_reg[62] , \edb_top_inst/la0/data_out_shift_reg[63] , 
        \edb_top_inst/la0/module_state[1] , \edb_top_inst/la0/module_state[2] , 
        \edb_top_inst/la0/module_state[3] , \edb_top_inst/la0/crc_data_out[0] , 
        \edb_top_inst/la0/crc_data_out[1] , \edb_top_inst/la0/crc_data_out[2] , 
        \edb_top_inst/la0/crc_data_out[3] , \edb_top_inst/la0/crc_data_out[4] , 
        \edb_top_inst/la0/crc_data_out[5] , \edb_top_inst/la0/crc_data_out[6] , 
        \edb_top_inst/la0/crc_data_out[7] , \edb_top_inst/la0/crc_data_out[8] , 
        \edb_top_inst/la0/crc_data_out[9] , \edb_top_inst/la0/crc_data_out[10] , 
        \edb_top_inst/la0/crc_data_out[11] , \edb_top_inst/la0/crc_data_out[12] , 
        \edb_top_inst/la0/crc_data_out[13] , \edb_top_inst/la0/crc_data_out[14] , 
        \edb_top_inst/la0/crc_data_out[15] , \edb_top_inst/la0/crc_data_out[16] , 
        \edb_top_inst/la0/crc_data_out[17] , \edb_top_inst/la0/crc_data_out[18] , 
        \edb_top_inst/la0/crc_data_out[19] , \edb_top_inst/la0/crc_data_out[20] , 
        \edb_top_inst/la0/crc_data_out[21] , \edb_top_inst/la0/crc_data_out[22] , 
        \edb_top_inst/la0/crc_data_out[23] , \edb_top_inst/la0/crc_data_out[24] , 
        \edb_top_inst/la0/crc_data_out[25] , \edb_top_inst/la0/crc_data_out[26] , 
        \edb_top_inst/la0/crc_data_out[27] , \edb_top_inst/la0/crc_data_out[28] , 
        \edb_top_inst/la0/crc_data_out[29] , \edb_top_inst/la0/crc_data_out[30] , 
        \edb_top_inst/la0/crc_data_out[31] , \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout , \edb_top_inst/la0/tu_trigger , 
        \edb_top_inst/la0/cap_fifo_din_cu[1] , \edb_top_inst/la0/cap_fifo_din_cu[2] , 
        \edb_top_inst/la0/cap_fifo_din_cu[5] , \edb_top_inst/la0/cap_fifo_din_cu[6] , 
        \edb_top_inst/la0/cap_fifo_din_cu[23] , \edb_top_inst/la0/cap_fifo_din_cu[40] , 
        \edb_top_inst/la0/cap_fifo_din_cu[41] , \edb_top_inst/la0/cap_fifo_din_tu[1] , 
        \edb_top_inst/la0/cap_fifo_din_tu[2] , \edb_top_inst/la0/cap_fifo_din_tu[5] , 
        \edb_top_inst/la0/cap_fifo_din_tu[6] , \edb_top_inst/la0/cap_fifo_din_tu[23] , 
        \edb_top_inst/la0/cap_fifo_din_tu[40] , \edb_top_inst/la0/cap_fifo_din_tu[41] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[0] , \edb_top_inst/la0/la_biu_inst/run_trig_p2 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , 
        \edb_top_inst/la0/la_biu_inst/str_sync , \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q , 
        \edb_top_inst/la0/data_from_biu[0] , \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[3] , \edb_top_inst/la0/la_biu_inst/curr_state[2] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[1] , \edb_top_inst/la0/biu_ready , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[15] , \edb_top_inst/la0/la_biu_inst/addr_reg[16] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[17] , \edb_top_inst/la0/la_biu_inst/addr_reg[18] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[19] , \edb_top_inst/la0/la_biu_inst/addr_reg[20] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[21] , \edb_top_inst/la0/la_biu_inst/addr_reg[22] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[23] , \edb_top_inst/la0/la_biu_inst/addr_reg[24] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[25] , \edb_top_inst/la0/la_biu_inst/addr_reg[26] , 
        \edb_top_inst/la0/data_from_biu[1] , \edb_top_inst/la0/data_from_biu[2] , 
        \edb_top_inst/la0/data_from_biu[3] , \edb_top_inst/la0/data_from_biu[4] , 
        \edb_top_inst/la0/data_from_biu[5] , \edb_top_inst/la0/data_from_biu[6] , 
        \edb_top_inst/la0/data_from_biu[7] , \edb_top_inst/la0/data_from_biu[8] , 
        \edb_top_inst/la0/data_from_biu[9] , \edb_top_inst/la0/data_from_biu[10] , 
        \edb_top_inst/la0/data_from_biu[11] , \edb_top_inst/la0/data_from_biu[12] , 
        \edb_top_inst/la0/data_from_biu[13] , \edb_top_inst/la0/data_from_biu[14] , 
        \edb_top_inst/la0/data_from_biu[15] , \edb_top_inst/la0/data_from_biu[16] , 
        \edb_top_inst/la0/data_from_biu[17] , \edb_top_inst/la0/data_from_biu[18] , 
        \edb_top_inst/la0/data_from_biu[19] , \edb_top_inst/la0/data_from_biu[20] , 
        \edb_top_inst/la0/data_from_biu[21] , \edb_top_inst/la0/data_from_biu[22] , 
        \edb_top_inst/la0/data_from_biu[23] , \edb_top_inst/la0/data_from_biu[24] , 
        \edb_top_inst/la0/data_from_biu[25] , \edb_top_inst/la0/data_from_biu[26] , 
        \edb_top_inst/la0/data_from_biu[27] , \edb_top_inst/la0/data_from_biu[28] , 
        \edb_top_inst/la0/data_from_biu[29] , \edb_top_inst/la0/data_from_biu[30] , 
        \edb_top_inst/la0/data_from_biu[31] , \edb_top_inst/la0/data_from_biu[32] , 
        \edb_top_inst/la0/data_from_biu[33] , \edb_top_inst/la0/data_from_biu[34] , 
        \edb_top_inst/la0/data_from_biu[35] , \edb_top_inst/la0/data_from_biu[36] , 
        \edb_top_inst/la0/data_from_biu[37] , \edb_top_inst/la0/data_from_biu[38] , 
        \edb_top_inst/la0/data_from_biu[39] , \edb_top_inst/la0/data_from_biu[40] , 
        \edb_top_inst/la0/data_from_biu[41] , \edb_top_inst/la0/data_from_biu[42] , 
        \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] , 
        \edb_top_inst/la0/la_sample_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[0] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] , 
        \edb_top_inst/la0/la_sample_cnt[1] , \edb_top_inst/la0/la_sample_cnt[2] , 
        \edb_top_inst/la0/la_sample_cnt[3] , \edb_top_inst/la0/la_sample_cnt[4] , 
        \edb_top_inst/la0/la_sample_cnt[5] , \edb_top_inst/la0/la_sample_cnt[6] , 
        \edb_top_inst/la0/la_sample_cnt[7] , \edb_top_inst/la0/la_sample_cnt[8] , 
        \edb_top_inst/la0/la_sample_cnt[9] , \edb_top_inst/la0/la_sample_cnt[10] , 
        \edb_top_inst/la0/la_sample_cnt[11] , \edb_top_inst/la0/la_sample_cnt[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[1] , \edb_top_inst/la0/la_biu_inst/fifo_counter[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[3] , \edb_top_inst/la0/la_biu_inst/fifo_counter[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[5] , \edb_top_inst/la0/la_biu_inst/fifo_counter[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[7] , \edb_top_inst/la0/la_biu_inst/fifo_counter[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[9] , \edb_top_inst/la0/la_biu_inst/fifo_counter[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[11] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] , 
        \edb_top_inst/la0/internal_register_select[1] , \edb_top_inst/la0/internal_register_select[2] , 
        \edb_top_inst/la0/internal_register_select[3] , \edb_top_inst/la0/internal_register_select[4] , 
        \edb_top_inst/la0/internal_register_select[5] , \edb_top_inst/la0/internal_register_select[6] , 
        \edb_top_inst/la0/internal_register_select[7] , \edb_top_inst/la0/internal_register_select[8] , 
        \edb_top_inst/la0/internal_register_select[9] , \edb_top_inst/la0/internal_register_select[10] , 
        \edb_top_inst/la0/internal_register_select[11] , \edb_top_inst/la0/internal_register_select[12] , 
        \edb_top_inst/la0/la_trig_pos[1] , \edb_top_inst/la0/la_trig_pos[2] , 
        \edb_top_inst/la0/la_trig_pos[3] , \edb_top_inst/la0/la_trig_pos[4] , 
        \edb_top_inst/la0/la_trig_pos[5] , \edb_top_inst/la0/la_trig_pos[6] , 
        \edb_top_inst/la0/la_trig_pos[7] , \edb_top_inst/la0/la_trig_pos[8] , 
        \edb_top_inst/la0/la_trig_pos[9] , \edb_top_inst/la0/la_trig_pos[10] , 
        \edb_top_inst/la0/la_trig_pos[11] , \edb_top_inst/la0/la_trig_pos[12] , 
        \edb_top_inst/la0/la_trig_pos[13] , \edb_top_inst/la0/la_trig_pos[14] , 
        \edb_top_inst/la0/la_trig_pos[15] , \edb_top_inst/la0/la_trig_pos[16] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[0] , \edb_top_inst/debug_hub_inst/module_id_reg[1] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[2] , \edb_top_inst/debug_hub_inst/module_id_reg[3] , 
        \edb_top_inst/n68 , \edb_top_inst/n70 , \edb_top_inst/n74 , \edb_top_inst/n694 , 
        \edb_top_inst/n696 , \edb_top_inst/n697 , \edb_top_inst/n698 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_pre , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre , 
        \edb_top_inst/n2760 , \edb_top_inst/n2761 , \edb_top_inst/n2762 , 
        \edb_top_inst/n2763 , \edb_top_inst/n2764 , \edb_top_inst/n2765 , 
        \edb_top_inst/n2766 , \edb_top_inst/n2767 , \edb_top_inst/n2768 , 
        \edb_top_inst/n2769 , \edb_top_inst/n2770 , \edb_top_inst/n2771 , 
        \edb_top_inst/n2772 , \edb_top_inst/n2773 , \edb_top_inst/n2774 , 
        \edb_top_inst/n2775 , \edb_top_inst/n2776 , \edb_top_inst/n2777 , 
        \edb_top_inst/n2778 , \edb_top_inst/n2779 , \edb_top_inst/n2780 , 
        \edb_top_inst/n2781 , \edb_top_inst/n2782 , \edb_top_inst/n2783 , 
        \edb_top_inst/n2784 , \edb_top_inst/n2785 , \edb_top_inst/n2786 , 
        \edb_top_inst/n2787 , \edb_top_inst/n2788 , \edb_top_inst/n2789 , 
        \edb_top_inst/n2790 , \edb_top_inst/n2791 , \edb_top_inst/n2792 , 
        \edb_top_inst/n2793 , \edb_top_inst/n2794 , \edb_top_inst/n2795 , 
        \edb_top_inst/n2796 , \edb_top_inst/n2797 , \edb_top_inst/n2798 , 
        \edb_top_inst/n2799 , \edb_top_inst/n2800 , \edb_top_inst/n2801 , 
        \edb_top_inst/n2802 , \edb_top_inst/n2803 , \edb_top_inst/n2804 , 
        \edb_top_inst/n2805 , \edb_top_inst/n2806 , \edb_top_inst/n2807 , 
        \edb_top_inst/n2808 , \edb_top_inst/n2809 , \edb_top_inst/n2810 , 
        \edb_top_inst/n2811 , \edb_top_inst/n2812 , \edb_top_inst/n2813 , 
        \edb_top_inst/n2814 , \edb_top_inst/n2815 , \edb_top_inst/n2816 , 
        \edb_top_inst/n2817 , \edb_top_inst/n2818 , \edb_top_inst/n2819 , 
        \edb_top_inst/n2820 , \edb_top_inst/n2736 , \edb_top_inst/n2733 , 
        \edb_top_inst/n2821 , \edb_top_inst/n1249 , \edb_top_inst/n2822 , 
        \edb_top_inst/n2823 , \edb_top_inst/n2824 , \edb_top_inst/n2825 , 
        \edb_top_inst/n2826 , \edb_top_inst/n2827 , \edb_top_inst/n2828 , 
        \edb_top_inst/n2829 , \edb_top_inst/n2830 , \edb_top_inst/n2831 , 
        \edb_top_inst/n2832 , \edb_top_inst/n2833 , \edb_top_inst/n2834 , 
        \edb_top_inst/n2835 , \edb_top_inst/n2836 , \edb_top_inst/n2837 , 
        \edb_top_inst/n2838 , \edb_top_inst/n2839 , \edb_top_inst/n2840 , 
        \edb_top_inst/n2841 , \edb_top_inst/n2842 , \edb_top_inst/n2843 , 
        \edb_top_inst/n2844 , \edb_top_inst/n2845 , \edb_top_inst/n2846 , 
        \edb_top_inst/n2847 , \edb_top_inst/n2848 , \edb_top_inst/n2849 , 
        \edb_top_inst/n2850 , \edb_top_inst/n2851 , \edb_top_inst/n2852 , 
        \edb_top_inst/n2853 , \edb_top_inst/n2854 , \edb_top_inst/n2855 , 
        \edb_top_inst/n2856 , \edb_top_inst/n2857 , \edb_top_inst/n2858 , 
        \edb_top_inst/n2859 , \edb_top_inst/n2860 , \edb_top_inst/n2861 , 
        \edb_top_inst/n2862 , \edb_top_inst/n2863 , \edb_top_inst/n2864 , 
        \edb_top_inst/n2865 , \edb_top_inst/n2866 , \edb_top_inst/n2867 , 
        \edb_top_inst/n2868 , \edb_top_inst/n2869 , \edb_top_inst/n2870 , 
        \edb_top_inst/n2871 , \edb_top_inst/n2872 , \edb_top_inst/n2873 , 
        \edb_top_inst/n2874 , \edb_top_inst/n2875 , \edb_top_inst/n2876 , 
        \edb_top_inst/n2877 , \edb_top_inst/n2878 , \edb_top_inst/n2879 , 
        \edb_top_inst/n2880 , \edb_top_inst/n2881 , \edb_top_inst/n2882 , 
        \edb_top_inst/n2888 , \edb_top_inst/n2889 , \edb_top_inst/n2890 , 
        \edb_top_inst/n2891 , \edb_top_inst/n2892 , \edb_top_inst/n2893 , 
        \edb_top_inst/n2894 , \edb_top_inst/n2895 , \edb_top_inst/n2896 , 
        \edb_top_inst/n2897 , \edb_top_inst/n2898 , \edb_top_inst/n2899 , 
        \edb_top_inst/n2900 , \edb_top_inst/n2901 , \edb_top_inst/n2902 , 
        \edb_top_inst/n2903 , \edb_top_inst/n2904 , \edb_top_inst/n2905 , 
        \edb_top_inst/n2906 , \edb_top_inst/n2907 , \edb_top_inst/n2908 , 
        \edb_top_inst/n2909 , \edb_top_inst/n2910 , \edb_top_inst/n2911 , 
        \edb_top_inst/n2912 , \edb_top_inst/n2913 , \edb_top_inst/n2914 , 
        \edb_top_inst/n2915 , \edb_top_inst/n2916 , \edb_top_inst/n2917 , 
        \edb_top_inst/n2918 , \edb_top_inst/n2919 , \edb_top_inst/n2920 , 
        \edb_top_inst/n2921 , \edb_top_inst/n2922 , \edb_top_inst/n2923 , 
        \edb_top_inst/n2924 , \edb_top_inst/n2925 , \edb_top_inst/n2926 , 
        \edb_top_inst/n2927 , \edb_top_inst/n2928 , \edb_top_inst/n2929 , 
        \edb_top_inst/n2930 , \edb_top_inst/n2931 , \edb_top_inst/n2932 , 
        \edb_top_inst/n2933 , \edb_top_inst/n2934 , \edb_top_inst/n2935 , 
        \edb_top_inst/n2936 , \edb_top_inst/n2937 , \edb_top_inst/n2938 , 
        \edb_top_inst/n2939 , \edb_top_inst/n2940 , \edb_top_inst/n2941 , 
        \edb_top_inst/n2942 , \edb_top_inst/n2943 , \edb_top_inst/n2944 , 
        \edb_top_inst/n2945 , \edb_top_inst/n2946 , \edb_top_inst/n2947 , 
        \edb_top_inst/n2948 , \edb_top_inst/n2949 , \edb_top_inst/n2950 , 
        \edb_top_inst/n2951 , \edb_top_inst/n2952 , \edb_top_inst/n2953 , 
        \edb_top_inst/n2954 , \edb_top_inst/n2955 , \edb_top_inst/n2956 , 
        \edb_top_inst/n2957 , \edb_top_inst/n2958 , \edb_top_inst/n2959 , 
        \edb_top_inst/n2960 , \edb_top_inst/n2961 , \edb_top_inst/n2962 , 
        \edb_top_inst/n2963 , \edb_top_inst/n2964 , \edb_top_inst/n2965 , 
        \edb_top_inst/n2966 , \edb_top_inst/n2967 , \edb_top_inst/n2968 , 
        \edb_top_inst/n2969 , \edb_top_inst/n2970 , \edb_top_inst/n2971 , 
        \edb_top_inst/n2972 , \edb_top_inst/n2973 , \edb_top_inst/n2974 , 
        \edb_top_inst/n2975 , \edb_top_inst/n2976 , \edb_top_inst/n2977 , 
        \edb_top_inst/n2978 , \edb_top_inst/n2979 , \edb_top_inst/n2980 , 
        \edb_top_inst/n2981 , \edb_top_inst/n2982 , \edb_top_inst/n2983 , 
        \edb_top_inst/n2984 , \edb_top_inst/n2985 , \edb_top_inst/n2986 , 
        \edb_top_inst/n2987 , \edb_top_inst/n2988 , \edb_top_inst/n2989 , 
        \edb_top_inst/n2990 , \edb_top_inst/n2991 , \edb_top_inst/n2992 , 
        \edb_top_inst/n2993 , \edb_top_inst/n2994 , \edb_top_inst/n2995 , 
        \edb_top_inst/n2996 , \edb_top_inst/n2997 , \edb_top_inst/n2998 , 
        \edb_top_inst/n2999 , \edb_top_inst/n3000 , \edb_top_inst/n3001 , 
        \edb_top_inst/n3002 , \edb_top_inst/n3003 , \edb_top_inst/n3004 , 
        \edb_top_inst/n3005 , \edb_top_inst/n3006 , \edb_top_inst/n3007 , 
        \edb_top_inst/n3008 , \edb_top_inst/n3009 , \edb_top_inst/n3010 , 
        \edb_top_inst/n3011 , \edb_top_inst/n3012 , \edb_top_inst/n3013 , 
        \edb_top_inst/n3014 , \edb_top_inst/n3015 , \edb_top_inst/n3016 , 
        \edb_top_inst/n3017 , \edb_top_inst/n3018 , \edb_top_inst/n3019 , 
        \edb_top_inst/n3020 , \edb_top_inst/n3021 , \edb_top_inst/n3022 , 
        \edb_top_inst/n3023 , \edb_top_inst/n3024 , \edb_top_inst/n3025 , 
        \edb_top_inst/n3026 , \edb_top_inst/n3027 , \edb_top_inst/n3028 , 
        \edb_top_inst/n3029 , \edb_top_inst/n3030 , \edb_top_inst/n3031 , 
        \edb_top_inst/n3032 , \edb_top_inst/n3033 , \edb_top_inst/n3034 , 
        \edb_top_inst/n3035 , \edb_top_inst/n3036 , \edb_top_inst/n3037 , 
        \edb_top_inst/n3038 , \edb_top_inst/n3039 , \edb_top_inst/n3040 , 
        \edb_top_inst/n3041 , \edb_top_inst/n3042 , \edb_top_inst/n3043 , 
        \edb_top_inst/n3044 , \edb_top_inst/n3045 , \edb_top_inst/n3046 , 
        \edb_top_inst/n3047 , \edb_top_inst/n3048 , \edb_top_inst/n3049 , 
        \edb_top_inst/n3050 , \edb_top_inst/n3051 , \edb_top_inst/n3052 , 
        \edb_top_inst/n3053 , \edb_top_inst/n3054 , \edb_top_inst/n3055 , 
        \edb_top_inst/n3056 , \edb_top_inst/n3057 , \edb_top_inst/n3058 , 
        \edb_top_inst/n3059 , \edb_top_inst/n3060 , \edb_top_inst/n3061 , 
        \edb_top_inst/n3062 , \edb_top_inst/n3063 , \edb_top_inst/n3064 , 
        \edb_top_inst/n3065 , \edb_top_inst/n3066 , \edb_top_inst/n3067 , 
        \edb_top_inst/n3068 , \edb_top_inst/n3069 , \edb_top_inst/n3070 , 
        \edb_top_inst/n3071 , \edb_top_inst/n3072 , \edb_top_inst/n3073 , 
        \edb_top_inst/n3074 , \edb_top_inst/n3075 , \edb_top_inst/n3076 , 
        \edb_top_inst/n3077 , \edb_top_inst/n3078 , \edb_top_inst/n3079 , 
        \edb_top_inst/n3080 , \edb_top_inst/n3081 , \edb_top_inst/n3082 , 
        \edb_top_inst/n3083 , \edb_top_inst/n3084 , \edb_top_inst/n3085 , 
        \edb_top_inst/n3086 , \edb_top_inst/n3087 , \edb_top_inst/n3088 , 
        \edb_top_inst/n3089 , \edb_top_inst/n3090 , \edb_top_inst/n3091 , 
        \edb_top_inst/n3092 , \edb_top_inst/n3093 , \edb_top_inst/n3094 , 
        \edb_top_inst/n3095 , \edb_top_inst/n3096 , \edb_top_inst/n3097 , 
        \edb_top_inst/n3098 , \edb_top_inst/n3099 , \edb_top_inst/n3100 , 
        \edb_top_inst/n3101 , \edb_top_inst/n3102 , \edb_top_inst/n3103 , 
        \edb_top_inst/n3104 , \edb_top_inst/n3105 , \edb_top_inst/n3106 , 
        \edb_top_inst/n3107 , \edb_top_inst/n3108 , \edb_top_inst/n3109 , 
        \edb_top_inst/n3110 , \edb_top_inst/n3111 , \edb_top_inst/n3112 , 
        \edb_top_inst/n3113 , \edb_top_inst/n3114 , \edb_top_inst/n3115 , 
        \edb_top_inst/n3116 , \edb_top_inst/n3117 , \edb_top_inst/n3118 , 
        \edb_top_inst/n3119 , \edb_top_inst/n3120 , \edb_top_inst/n3121 , 
        \edb_top_inst/n3122 , \edb_top_inst/n3123 , \edb_top_inst/n3124 , 
        \edb_top_inst/n3125 , \edb_top_inst/n3126 , \edb_top_inst/n3127 , 
        \edb_top_inst/n3128 , \edb_top_inst/n3129 , \edb_top_inst/n3130 , 
        \edb_top_inst/n3131 , \edb_top_inst/n3132 , \edb_top_inst/n3133 , 
        \edb_top_inst/n3134 , \edb_top_inst/n3135 , \edb_top_inst/n3136 , 
        \edb_top_inst/n3137 , \edb_top_inst/n3138 , \edb_top_inst/n3139 , 
        \edb_top_inst/n3140 , \edb_top_inst/n3141 , \edb_top_inst/n3142 , 
        \edb_top_inst/n3143 , \edb_top_inst/n3144 , \edb_top_inst/n3145 , 
        \edb_top_inst/n3146 , \edb_top_inst/n3147 , \edb_top_inst/n3148 , 
        \edb_top_inst/n3149 , \edb_top_inst/n3150 , \edb_top_inst/n3151 , 
        \edb_top_inst/n3152 , \edb_top_inst/n3153 , \edb_top_inst/n3154 , 
        \edb_top_inst/n3155 , \edb_top_inst/n3156 , \edb_top_inst/n3157 , 
        \edb_top_inst/n3158 , \edb_top_inst/n3159 , \edb_top_inst/n3160 , 
        \edb_top_inst/n3161 , \edb_top_inst/n3162 , \edb_top_inst/n3163 , 
        \edb_top_inst/n3164 , \edb_top_inst/n3165 , \edb_top_inst/n3166 , 
        \edb_top_inst/n3167 , \edb_top_inst/n3168 , \edb_top_inst/n3169 , 
        \edb_top_inst/n3170 , \edb_top_inst/n3171 , \edb_top_inst/n3172 , 
        \edb_top_inst/n3173 , \edb_top_inst/n3174 , \edb_top_inst/n3175 , 
        \edb_top_inst/n3176 , \edb_top_inst/n3177 , \edb_top_inst/n3178 , 
        \edb_top_inst/n3179 , \edb_top_inst/n3180 , \edb_top_inst/n3181 , 
        \edb_top_inst/n3182 , \edb_top_inst/n3183 , \edb_top_inst/n3184 , 
        \edb_top_inst/n3185 , \edb_top_inst/n3186 , \edb_top_inst/n3187 , 
        \edb_top_inst/n3188 , \edb_top_inst/n3189 , \edb_top_inst/n3190 , 
        \edb_top_inst/n3191 , \edb_top_inst/n3192 , \edb_top_inst/n3193 , 
        \edb_top_inst/n3194 , \edb_top_inst/n3195 , \edb_top_inst/n3196 , 
        \edb_top_inst/n3197 , \edb_top_inst/n3198 , \edb_top_inst/n3199 , 
        \edb_top_inst/n3200 , \edb_top_inst/n3201 , \edb_top_inst/n3202 , 
        \edb_top_inst/n3203 , \edb_top_inst/n3204 , \edb_top_inst/n3205 , 
        \edb_top_inst/n3206 , \edb_top_inst/n3207 , \edb_top_inst/n3208 , 
        \edb_top_inst/n3209 , \edb_top_inst/n3210 , \edb_top_inst/n3211 , 
        \edb_top_inst/n3212 , \edb_top_inst/n3213 , \edb_top_inst/n3214 , 
        \edb_top_inst/n3215 , \edb_top_inst/n3216 , \edb_top_inst/n3217 , 
        \edb_top_inst/n3218 , \edb_top_inst/n3219 , \edb_top_inst/n3220 , 
        \edb_top_inst/n3221 , \edb_top_inst/n3222 , \edb_top_inst/n3223 , 
        \edb_top_inst/n3224 , \edb_top_inst/n3225 , \edb_top_inst/n3226 , 
        \edb_top_inst/n3227 , \edb_top_inst/n3228 , \edb_top_inst/n3229 , 
        \edb_top_inst/n3230 , \edb_top_inst/n3231 , \edb_top_inst/n3232 , 
        \edb_top_inst/n3233 , \edb_top_inst/n3234 , \edb_top_inst/n3235 , 
        \edb_top_inst/n3236 , \edb_top_inst/n3237 , \edb_top_inst/n3238 , 
        \edb_top_inst/n3239 , \edb_top_inst/n3240 , \edb_top_inst/n3241 , 
        \edb_top_inst/n3242 , \edb_top_inst/n3243 , \edb_top_inst/n3244 , 
        \edb_top_inst/n3245 , \edb_top_inst/n3246 , \edb_top_inst/n3247 , 
        \edb_top_inst/n3248 , \edb_top_inst/n3249 , \edb_top_inst/n3250 , 
        \edb_top_inst/n3251 , \edb_top_inst/n3252 , \edb_top_inst/n3253 , 
        \edb_top_inst/n3254 , \edb_top_inst/n3255 , \edb_top_inst/n3256 , 
        \edb_top_inst/n3257 , \edb_top_inst/n3258 , \edb_top_inst/n3259 , 
        \edb_top_inst/n3260 , \edb_top_inst/n3261 , \edb_top_inst/n3262 , 
        \edb_top_inst/n3263 , \edb_top_inst/n3264 , \edb_top_inst/n3265 , 
        \edb_top_inst/n3266 , \edb_top_inst/n3267 , \edb_top_inst/n3268 , 
        \edb_top_inst/n3269 , \edb_top_inst/n3270 , \edb_top_inst/n3271 , 
        \edb_top_inst/n3272 , \edb_top_inst/n3273 , \edb_top_inst/n3274 , 
        \edb_top_inst/n3275 , \edb_top_inst/n3276 , \edb_top_inst/n3277 , 
        \edb_top_inst/n3278 , \edb_top_inst/n3279 , \edb_top_inst/n3280 , 
        \edb_top_inst/n3281 , \edb_top_inst/n3282 , \edb_top_inst/n3283 , 
        \edb_top_inst/n3284 , \edb_top_inst/n3285 , \edb_top_inst/n3286 , 
        \edb_top_inst/n3287 , \edb_top_inst/n3288 , \edb_top_inst/n3289 , 
        \edb_top_inst/n3290 , \edb_top_inst/n3291 , \edb_top_inst/n3292 , 
        \edb_top_inst/n3293 , \edb_top_inst/n3294 , \edb_top_inst/n3295 , 
        \edb_top_inst/n3296 , \edb_top_inst/n3297 , \edb_top_inst/n3298 , 
        \edb_top_inst/n3299 , \edb_top_inst/n3300 , \edb_top_inst/n3301 , 
        \edb_top_inst/n3302 , \edb_top_inst/n3303 , \edb_top_inst/n3304 , 
        \edb_top_inst/n3305 , \edb_top_inst/n3306 , \edb_top_inst/n3307 , 
        \edb_top_inst/n3308 , \edb_top_inst/n3309 , \edb_top_inst/n3310 , 
        \edb_top_inst/n3311 , \edb_top_inst/n3312 , \edb_top_inst/n3313 , 
        \edb_top_inst/n3314 , \edb_top_inst/n3315 , \edb_top_inst/n3316 , 
        \edb_top_inst/n3317 , \edb_top_inst/n3318 , \edb_top_inst/n3319 , 
        \edb_top_inst/n3320 , \edb_top_inst/n3321 , \edb_top_inst/n3322 , 
        \edb_top_inst/n3323 , \edb_top_inst/n3324 , \edb_top_inst/n3325 , 
        \edb_top_inst/n3326 , \edb_top_inst/n3327 , \edb_top_inst/n3328 , 
        \edb_top_inst/n3329 , \edb_top_inst/n3330 , \edb_top_inst/n3331 , 
        \edb_top_inst/n3332 , \edb_top_inst/n3333 , \edb_top_inst/n3334 , 
        \edb_top_inst/n3335 , \edb_top_inst/n3336 , \edb_top_inst/n3337 , 
        \edb_top_inst/n3338 , \edb_top_inst/n3339 , \edb_top_inst/n3340 , 
        \edb_top_inst/n2739 , \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0 , 
        \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 , n2823, n2824, 
        n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
        n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, 
        n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, 
        n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, 
        n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, 
        n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, 
        n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, 
        n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, 
        n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, 
        n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, 
        n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, 
        n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
        n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
        n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, 
        n2937, n2938, n2946, n2947, n2948, n2949, n2950, n2951, 
        n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, 
        n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, 
        n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, 
        n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
        n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, 
        n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
        n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, 
        n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, 
        n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
        n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, 
        n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, 
        n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, 
        n3048, n3049, wCdcFifoFull, rSRST, \MCsiRxController/n281 , 
        \MCsiRxController/MCsi2Decoder/n631 , \MCsiRxController/MCsi2Decoder/n633 , 
        \MCsiRxController/MCsi2Decoder/n7 , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[0] , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qFullAllmost , 
        \MCsiRxController/MCsi2Decoder/n585 , \MCsiRxController/MCsi2Decoder/n604 , 
        \MCsiRxController/MCsi2Decoder/qLineCntRst , \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE , 
        \MCsiRxController/MCsi2Decoder/n97 , \MCsiRxController/MCsi2Decoder/n607 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n19 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n233 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n238 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n243 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n248 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n253 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n258 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n263 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n268 , 
        \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n273 , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] , 
        \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[1] , \MCsiRxController/MCsi2Decoder/wFtiRd[2] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[3] , \MCsiRxController/MCsi2Decoder/wFtiRd[4] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[5] , \MCsiRxController/MCsi2Decoder/wFtiRd[6] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[7] , \MCsiRxController/MCsi2Decoder/wFtiRd[8] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[9] , \MCsiRxController/MCsi2Decoder/wFtiRd[10] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[11] , \MCsiRxController/MCsi2Decoder/wFtiRd[12] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[13] , \MCsiRxController/MCsi2Decoder/wFtiRd[14] , 
        \MCsiRxController/MCsi2Decoder/wFtiRd[15] , \MCsiRxController/MCsi2Decoder/equal_63/n5 , 
        \MCsiRxController/MCsi2Decoder/equal_60/n5 , \MCsiRxController/genblk1[0].mVideoFIFO/qRE , 
        \MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost , \MCsiRxController/genblk1[0].mVideoFIFO/qRVD , 
        \MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 , \MCsiRxController/genblk1[0].mVideoFIFO/n436 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n441 , \MCsiRxController/genblk1[0].mVideoFIFO/n446 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n451 , \MCsiRxController/genblk1[0].mVideoFIFO/n456 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n461 , \MCsiRxController/genblk1[0].mVideoFIFO/n466 , 
        \MCsiRxController/genblk1[0].mVideoFIFO/n471 , \MCsiRxController/n280 , 
        \MCsiRxController/n279 , \MCsiRxController/n278 , \MCsiRxController/n277 , 
        \MCsiRxController/n276 , \MCsiRxController/n275 , \MCsiRxController/n274 , 
        \MCsiRxController/n273 , \MCsiRxController/n272 , \MCsiRxController/n271 , 
        \MCsiRxController/n270 , \MCsiRxController/n269 , \MCsiRxController/n268 , 
        \MCsiRxController/n267 , \MCsiRxController/n266 , \MVideoPostProcess/qVtgRstCntCke , 
        \MVideoPostProcess/rVtgRstSel , \MVideoPostProcess/equal_18/n21 , 
        \~n1835 , ceg_net939, \MVideoPostProcess/inst_adv7511_config/n816 , 
        \MVideoPostProcess/inst_adv7511_config/n833 , \~ceg_net512 , \MVideoPostProcess/inst_adv7511_config/n268 , 
        ceg_net995, \MVideoPostProcess/inst_adv7511_config/n1107 , \MVideoPostProcess/inst_adv7511_config/n1224 , 
        \MVideoPostProcess/inst_adv7511_config/n277 , ceg_net479, ceg_net43, 
        ceg_net1327, \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] , 
        \MVideoPostProcess/inst_adv7511_config/n1243 , \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 , 
        ceg_net1087, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 , 
        ceg_net1335, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 , 
        ceg_net566, \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] , 
        ceg_net1400, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 , 
        ceg_net1463, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 , 
        ceg_net1361, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 , 
        ceg_net616, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 , 
        \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 , 
        ceg_net1471, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 , 
        ceg_net1480, \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 , 
        ceg_net1488, n8455, n8454, n8453, n8452, \MVideoPostProcess/mVideoTimingGen/qVrange , 
        \MVideoPostProcess/inst_adv7511_config/n251 , \MVideoPostProcess/inst_adv7511_config/n250 , 
        \MVideoPostProcess/inst_adv7511_config/n249 , \MVideoPostProcess/inst_adv7511_config/n248 , 
        \MVideoPostProcess/inst_adv7511_config/n247 , \MVideoPostProcess/inst_adv7511_config/n246 , 
        \MVideoPostProcess/inst_adv7511_config/n245 , \MVideoPostProcess/inst_adv7511_config/n244 , 
        \MVideoPostProcess/inst_adv7511_config/n700 , \MVideoPostProcess/inst_adv7511_config/n705 , 
        \MVideoPostProcess/inst_adv7511_config/n710 , \MVideoPostProcess/inst_adv7511_config/n715 , 
        \MVideoPostProcess/inst_adv7511_config/n720 , \MVideoPostProcess/inst_adv7511_config/n725 , 
        \MVideoPostProcess/inst_adv7511_config/n730 , \MVideoPostProcess/inst_adv7511_config/n735 , 
        \MVideoPostProcess/inst_adv7511_config/n740 , \MVideoPostProcess/inst_adv7511_config/n745 , 
        \MVideoPostProcess/inst_adv7511_config/n750 , \MVideoPostProcess/inst_adv7511_config/n755 , 
        \MVideoPostProcess/inst_adv7511_config/n760 , \MVideoPostProcess/inst_adv7511_config/n765 , 
        \MVideoPostProcess/inst_adv7511_config/n770 , \MVideoPostProcess/inst_adv7511_config/n780 , 
        \MVideoPostProcess/inst_adv7511_config/n785 , \MVideoPostProcess/inst_adv7511_config/n790 , 
        \MVideoPostProcess/inst_adv7511_config/n795 , \MVideoPostProcess/inst_adv7511_config/n800 , 
        \MVideoPostProcess/inst_adv7511_config/n805 , \MVideoPostProcess/inst_adv7511_config/n810 , 
        \MVideoPostProcess/inst_adv7511_config/n276 , \MVideoPostProcess/inst_adv7511_config/n275 , 
        \MVideoPostProcess/inst_adv7511_config/n274 , \MVideoPostProcess/inst_adv7511_config/n273 , 
        \MVideoPostProcess/inst_adv7511_config/n272 , \MVideoPostProcess/inst_adv7511_config/n271 , 
        \MVideoPostProcess/inst_adv7511_config/n270 , \MVideoPostProcess/mVideoTimingGen/n131 , 
        \MVideoPostProcess/mVideoTimingGen/equal_12/n23 , \MVideoPostProcess/rVtgRST[2] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] , 
        \MVideoPostProcess/mVideoTimingGen/qVde , \MVideoPostProcess/mVideoTimingGen/n267 , 
        \MVideoPostProcess/mVideoTimingGen/rHSync[3] , \MVideoPostProcess/mVideoTimingGen/n130 , 
        \MVideoPostProcess/mVideoTimingGen/n129 , \MVideoPostProcess/mVideoTimingGen/n126 , 
        \MVideoPostProcess/mVideoTimingGen/n125 , \MVideoPostProcess/mVideoTimingGen/n121 , 
        \MVideoPostProcess/mVideoTimingGen/qHrange , \MVideoPostProcess/mVideoTimingGen/rVSync[3] , 
        \MVideoPostProcess/wVgaGenFDe , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n433 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n438 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n443 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n448 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n453 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n458 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n463 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n468 , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n473 , 
        \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] , 
        \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] , 
        \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] , 
        \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] , 
        \genblk1.genblk1[0].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[0].mPulseGenerator/equal_12/n23 , 
        \genblk1.genblk1[1].mPulseGenerator/equal_6/n5 , \genblk1.genblk1[1].mPulseGenerator/equal_12/n3 , 
        \genblk1.genblk1[1].mPulseGenerator/n50 , \genblk1.genblk1[3].mPulseGenerator/equal_6/n5 , 
        \genblk1.genblk1[3].mPulseGenerator/n50 , \genblk1.genblk1[4].mPulseGenerator/equal_6/n5 , 
        \genblk1.genblk1[4].mPulseGenerator/n50 , \edb_top_inst/la0/n1340 , 
        \edb_top_inst/ceg_net5 , \edb_top_inst/edb_user_dr[60] , \edb_top_inst/la0/n1312 , 
        \edb_top_inst/la0/n1341 , \edb_top_inst/la0/n1342 , \edb_top_inst/edb_user_dr[62] , 
        \edb_top_inst/edb_user_dr[0] , \edb_top_inst/la0/n1396 , \edb_top_inst/edb_user_dr[42] , 
        \edb_top_inst/la0/n1913 , \edb_top_inst/edb_user_dr[59] , \edb_top_inst/la0/n1965 , 
        \edb_top_inst/la0/data_to_addr_counter[0] , \edb_top_inst/la0/addr_ct_en , 
        \edb_top_inst/edb_user_dr[77] , \edb_top_inst/la0/op_reg_en , \edb_top_inst/la0/n2189 , 
        \edb_top_inst/ceg_net26 , \edb_top_inst/la0/data_to_word_counter[0] , 
        \edb_top_inst/la0/word_ct_en , \edb_top_inst/la0/n2466 , \edb_top_inst/ceg_net14 , 
        \edb_top_inst/la0/module_next_state[0] , la0_probe1, \edb_top_inst/la0/n5294 , 
        \edb_top_inst/la0/n5492 , \edb_top_inst/la0/n6947 , \edb_top_inst/la0/n7907 , 
        \edb_top_inst/la0/n8105 , \edb_top_inst/la0/n8741 , \edb_top_inst/la0/n9645 , 
        \edb_top_inst/la0/n9843 , \edb_top_inst/la0/n10527 , \edb_top_inst/la0/n10542 , 
        \edb_top_inst/la0/n10740 , \edb_top_inst/la0/n11368 , \edb_top_inst/la0/n12201 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/edb_user_dr[64] , \edb_top_inst/la0/regsel_ld_en , 
        \edb_top_inst/edb_user_dr[43] , \edb_top_inst/edb_user_dr[61] , 
        \edb_top_inst/edb_user_dr[63] , \edb_top_inst/edb_user_dr[1] , \edb_top_inst/edb_user_dr[2] , 
        \edb_top_inst/edb_user_dr[3] , \edb_top_inst/edb_user_dr[4] , \edb_top_inst/edb_user_dr[5] , 
        \edb_top_inst/edb_user_dr[6] , \edb_top_inst/edb_user_dr[7] , \edb_top_inst/edb_user_dr[8] , 
        \edb_top_inst/edb_user_dr[9] , \edb_top_inst/edb_user_dr[10] , \edb_top_inst/edb_user_dr[11] , 
        \edb_top_inst/edb_user_dr[12] , \edb_top_inst/edb_user_dr[13] , 
        \edb_top_inst/edb_user_dr[14] , \edb_top_inst/edb_user_dr[15] , 
        \edb_top_inst/edb_user_dr[16] , \edb_top_inst/edb_user_dr[17] , 
        \edb_top_inst/edb_user_dr[18] , \edb_top_inst/edb_user_dr[19] , 
        \edb_top_inst/edb_user_dr[20] , \edb_top_inst/edb_user_dr[21] , 
        \edb_top_inst/edb_user_dr[22] , \edb_top_inst/edb_user_dr[23] , 
        \edb_top_inst/edb_user_dr[24] , \edb_top_inst/edb_user_dr[25] , 
        \edb_top_inst/edb_user_dr[26] , \edb_top_inst/edb_user_dr[27] , 
        \edb_top_inst/edb_user_dr[28] , \edb_top_inst/edb_user_dr[29] , 
        \edb_top_inst/edb_user_dr[30] , \edb_top_inst/edb_user_dr[31] , 
        \edb_top_inst/edb_user_dr[32] , \edb_top_inst/edb_user_dr[33] , 
        \edb_top_inst/edb_user_dr[34] , \edb_top_inst/edb_user_dr[35] , 
        \edb_top_inst/edb_user_dr[36] , \edb_top_inst/edb_user_dr[37] , 
        \edb_top_inst/edb_user_dr[38] , \edb_top_inst/edb_user_dr[39] , 
        \edb_top_inst/edb_user_dr[40] , \edb_top_inst/edb_user_dr[41] , 
        \edb_top_inst/edb_user_dr[44] , \edb_top_inst/edb_user_dr[45] , 
        \edb_top_inst/edb_user_dr[46] , \edb_top_inst/edb_user_dr[47] , 
        \edb_top_inst/edb_user_dr[48] , \edb_top_inst/edb_user_dr[49] , 
        \edb_top_inst/edb_user_dr[50] , \edb_top_inst/edb_user_dr[51] , 
        \edb_top_inst/edb_user_dr[52] , \edb_top_inst/edb_user_dr[53] , 
        \edb_top_inst/edb_user_dr[54] , \edb_top_inst/edb_user_dr[55] , 
        \edb_top_inst/edb_user_dr[56] , \edb_top_inst/edb_user_dr[57] , 
        \edb_top_inst/edb_user_dr[58] , \edb_top_inst/la0/data_to_addr_counter[1] , 
        \edb_top_inst/la0/data_to_addr_counter[2] , \edb_top_inst/la0/data_to_addr_counter[3] , 
        \edb_top_inst/la0/data_to_addr_counter[4] , \edb_top_inst/la0/data_to_addr_counter[5] , 
        \edb_top_inst/la0/data_to_addr_counter[6] , \edb_top_inst/la0/data_to_addr_counter[7] , 
        \edb_top_inst/la0/data_to_addr_counter[8] , \edb_top_inst/la0/data_to_addr_counter[9] , 
        \edb_top_inst/la0/data_to_addr_counter[10] , \edb_top_inst/la0/data_to_addr_counter[11] , 
        \edb_top_inst/la0/data_to_addr_counter[12] , \edb_top_inst/la0/data_to_addr_counter[13] , 
        \edb_top_inst/la0/data_to_addr_counter[14] , \edb_top_inst/la0/data_to_addr_counter[15] , 
        \edb_top_inst/la0/data_to_addr_counter[16] , \edb_top_inst/la0/data_to_addr_counter[17] , 
        \edb_top_inst/la0/data_to_addr_counter[18] , \edb_top_inst/la0/data_to_addr_counter[19] , 
        \edb_top_inst/la0/data_to_addr_counter[20] , \edb_top_inst/la0/data_to_addr_counter[21] , 
        \edb_top_inst/la0/data_to_addr_counter[22] , \edb_top_inst/la0/data_to_addr_counter[23] , 
        \edb_top_inst/la0/data_to_addr_counter[24] , \edb_top_inst/la0/data_to_addr_counter[25] , 
        \edb_top_inst/la0/data_to_addr_counter[26] , \edb_top_inst/edb_user_dr[78] , 
        \edb_top_inst/edb_user_dr[79] , \edb_top_inst/edb_user_dr[80] , 
        \edb_top_inst/la0/n2188 , \edb_top_inst/la0/n2187 , \edb_top_inst/la0/n2186 , 
        \edb_top_inst/la0/n2185 , \edb_top_inst/la0/n2184 , \edb_top_inst/la0/data_to_word_counter[1] , 
        \edb_top_inst/la0/data_to_word_counter[2] , \edb_top_inst/la0/data_to_word_counter[3] , 
        \edb_top_inst/la0/data_to_word_counter[4] , \edb_top_inst/la0/data_to_word_counter[5] , 
        \edb_top_inst/la0/data_to_word_counter[6] , \edb_top_inst/la0/data_to_word_counter[7] , 
        \edb_top_inst/la0/data_to_word_counter[8] , \edb_top_inst/la0/data_to_word_counter[9] , 
        \edb_top_inst/la0/data_to_word_counter[10] , \edb_top_inst/la0/data_to_word_counter[11] , 
        \edb_top_inst/la0/data_to_word_counter[12] , \edb_top_inst/la0/data_to_word_counter[13] , 
        \edb_top_inst/la0/data_to_word_counter[14] , \edb_top_inst/la0/data_to_word_counter[15] , 
        \edb_top_inst/la0/n2465 , \edb_top_inst/la0/n2464 , \edb_top_inst/la0/n2463 , 
        \edb_top_inst/la0/n2462 , \edb_top_inst/la0/n2461 , \edb_top_inst/la0/n2460 , 
        \edb_top_inst/la0/n2459 , \edb_top_inst/la0/n2458 , \edb_top_inst/la0/n2457 , 
        \edb_top_inst/la0/n2456 , \edb_top_inst/la0/n2455 , \edb_top_inst/la0/n2454 , 
        \edb_top_inst/la0/n2453 , \edb_top_inst/la0/n2452 , \edb_top_inst/la0/n2451 , 
        \edb_top_inst/la0/n2450 , \edb_top_inst/la0/n2449 , \edb_top_inst/la0/n2448 , 
        \edb_top_inst/la0/n2447 , \edb_top_inst/la0/n2446 , \edb_top_inst/la0/n2445 , 
        \edb_top_inst/la0/n2444 , \edb_top_inst/la0/n2443 , \edb_top_inst/la0/n2442 , 
        \edb_top_inst/la0/n2441 , \edb_top_inst/la0/n2440 , \edb_top_inst/la0/n2439 , 
        \edb_top_inst/la0/n2438 , \edb_top_inst/la0/n2437 , \edb_top_inst/la0/n2436 , 
        \edb_top_inst/la0/n2435 , \edb_top_inst/la0/n2434 , \edb_top_inst/la0/n2433 , 
        \edb_top_inst/la0/n2432 , \edb_top_inst/la0/n2431 , \edb_top_inst/la0/n2430 , 
        \edb_top_inst/la0/n2429 , \edb_top_inst/la0/n2428 , \edb_top_inst/la0/n2427 , 
        \edb_top_inst/la0/n2426 , \edb_top_inst/la0/n2425 , \edb_top_inst/la0/n2424 , 
        \edb_top_inst/la0/n2423 , \edb_top_inst/la0/n2422 , \edb_top_inst/la0/n2421 , 
        \edb_top_inst/la0/n2420 , \edb_top_inst/la0/n2419 , \edb_top_inst/la0/n2418 , 
        \edb_top_inst/la0/n2417 , \edb_top_inst/la0/n2416 , \edb_top_inst/la0/n2415 , 
        \edb_top_inst/la0/n2414 , \edb_top_inst/la0/n2413 , \edb_top_inst/la0/n2412 , 
        \edb_top_inst/la0/n2411 , \edb_top_inst/la0/n2410 , \edb_top_inst/la0/n2409 , 
        \edb_top_inst/la0/n2408 , \edb_top_inst/la0/n2407 , \edb_top_inst/la0/n2406 , 
        \edb_top_inst/la0/n2405 , \edb_top_inst/la0/n2404 , \edb_top_inst/la0/n2403 , 
        \edb_top_inst/la0/module_next_state[1] , \edb_top_inst/la0/module_next_state[2] , 
        \edb_top_inst/la0/module_next_state[3] , \edb_top_inst/la0/axi_crc_i/n150 , 
        \edb_top_inst/ceg_net221 , \edb_top_inst/la0/axi_crc_i/n149 , \edb_top_inst/la0/axi_crc_i/n148 , 
        \edb_top_inst/la0/axi_crc_i/n147 , \edb_top_inst/la0/axi_crc_i/n146 , 
        \edb_top_inst/la0/axi_crc_i/n145 , \edb_top_inst/la0/axi_crc_i/n144 , 
        \edb_top_inst/la0/axi_crc_i/n143 , \edb_top_inst/la0/axi_crc_i/n142 , 
        \edb_top_inst/la0/axi_crc_i/n141 , \edb_top_inst/la0/axi_crc_i/n140 , 
        \edb_top_inst/la0/axi_crc_i/n139 , \edb_top_inst/la0/axi_crc_i/n138 , 
        \edb_top_inst/la0/axi_crc_i/n137 , \edb_top_inst/la0/axi_crc_i/n136 , 
        \edb_top_inst/la0/axi_crc_i/n135 , \edb_top_inst/la0/axi_crc_i/n134 , 
        \edb_top_inst/la0/axi_crc_i/n133 , \edb_top_inst/la0/axi_crc_i/n132 , 
        \edb_top_inst/la0/axi_crc_i/n131 , \edb_top_inst/la0/axi_crc_i/n130 , 
        \edb_top_inst/la0/axi_crc_i/n129 , \edb_top_inst/la0/axi_crc_i/n128 , 
        \edb_top_inst/la0/axi_crc_i/n127 , \edb_top_inst/la0/axi_crc_i/n126 , 
        \edb_top_inst/la0/axi_crc_i/n125 , \edb_top_inst/la0/axi_crc_i/n124 , 
        \edb_top_inst/la0/axi_crc_i/n123 , \edb_top_inst/la0/axi_crc_i/n122 , 
        \edb_top_inst/la0/axi_crc_i/n121 , \edb_top_inst/la0/axi_crc_i/n120 , 
        \edb_top_inst/la0/axi_crc_i/n119 , \edb_top_inst/la0/n2766 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n3599 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n4432 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n5279 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n16 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n10 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n3 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n15 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n9 , \edb_top_inst/la0/n6114 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n7892 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n72 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n73 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n31 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n82 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n71 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n32 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n31 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n30 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n29 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n28 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n27 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n26 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n25 , \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n24 , 
        \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/n9630 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n38 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n36 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n34 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n21 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n15 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n38 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n36 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n21 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n15 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 , \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/trigger_tu/n89 , 
        \edb_top_inst/la0/la_biu_inst/next_state[0] , \edb_top_inst/la0/la_biu_inst/run_trig_p1 , 
        \edb_top_inst/la0/la_biu_inst/n382 , \edb_top_inst/la0/la_biu_inst/n1315 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[0] , \edb_top_inst/la0/la_biu_inst/next_fsm_state[0] , 
        \edb_top_inst/ceg_net351 , \edb_top_inst/la0/la_biu_inst/n1300 , 
        \edb_top_inst/la0/n17781 , \edb_top_inst/la0/la_biu_inst/next_state[2] , 
        \edb_top_inst/la0/la_biu_inst/next_state[1] , \edb_top_inst/ceg_net348 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[3] , \edb_top_inst/la0/la_biu_inst/fifo_dout[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[5] , \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[7] , \edb_top_inst/la0/la_biu_inst/fifo_dout[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[9] , \edb_top_inst/la0/la_biu_inst/fifo_dout[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[11] , \edb_top_inst/la0/la_biu_inst/fifo_dout[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[13] , \edb_top_inst/la0/la_biu_inst/fifo_dout[14] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[15] , \edb_top_inst/la0/la_biu_inst/fifo_dout[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[17] , \edb_top_inst/la0/la_biu_inst/fifo_dout[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[19] , \edb_top_inst/la0/la_biu_inst/fifo_dout[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[21] , \edb_top_inst/la0/la_biu_inst/fifo_dout[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[23] , \edb_top_inst/la0/la_biu_inst/fifo_dout[24] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[25] , \edb_top_inst/la0/la_biu_inst/fifo_dout[26] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[27] , \edb_top_inst/la0/la_biu_inst/fifo_dout[28] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[29] , \edb_top_inst/la0/la_biu_inst/fifo_dout[30] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[31] , \edb_top_inst/la0/la_biu_inst/fifo_dout[32] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[33] , \edb_top_inst/la0/la_biu_inst/fifo_dout[34] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[35] , \edb_top_inst/la0/la_biu_inst/fifo_dout[36] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[37] , \edb_top_inst/la0/la_biu_inst/fifo_dout[38] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[39] , \edb_top_inst/la0/la_biu_inst/fifo_dout[40] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[41] , \edb_top_inst/la0/la_biu_inst/fifo_dout[42] , 
        \edb_top_inst/la0/la_biu_inst/next_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , 
        \edb_top_inst/la0/la_biu_inst/fifo_rstn , \edb_top_inst/la0/la_biu_inst/n2053 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 , \edb_top_inst/la0/la_biu_inst/fifo_push , 
        \edb_top_inst/ceg_net355 , \edb_top_inst/n73 , \edb_top_inst/n1044 , 
        \edb_top_inst/n1042 , \edb_top_inst/n1040 , \edb_top_inst/n1038 , 
        \edb_top_inst/n1036 , \edb_top_inst/n1034 , \edb_top_inst/n1032 , 
        \edb_top_inst/n1030 , \edb_top_inst/n1028 , \edb_top_inst/n1027 , 
        \edb_top_inst/n693 , \edb_top_inst/n1025 , \edb_top_inst/n1023 , 
        \edb_top_inst/n1021 , \edb_top_inst/n1019 , \edb_top_inst/n1017 , 
        \edb_top_inst/n1015 , \edb_top_inst/n1013 , \edb_top_inst/n1011 , 
        \edb_top_inst/n1008 , \edb_top_inst/n1005 , \edb_top_inst/n695 , 
        \edb_top_inst/n856 , \edb_top_inst/n854 , \edb_top_inst/n852 , 
        \edb_top_inst/n850 , \edb_top_inst/n848 , \edb_top_inst/n846 , 
        \edb_top_inst/n844 , \edb_top_inst/n842 , \edb_top_inst/n840 , 
        \edb_top_inst/n838 , \edb_top_inst/n710 , \edb_top_inst/n731 , 
        \edb_top_inst/n729 , \edb_top_inst/n727 , \edb_top_inst/n725 , 
        \edb_top_inst/n723 , \edb_top_inst/n721 , \edb_top_inst/n719 , 
        \edb_top_inst/n717 , \edb_top_inst/n715 , \edb_top_inst/n713 , 
        \edb_top_inst/n712 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] , 
        \edb_top_inst/n711 , \edb_top_inst/n752 , \edb_top_inst/n750 , 
        \edb_top_inst/n748 , \edb_top_inst/n746 , \edb_top_inst/n744 , 
        \edb_top_inst/n742 , \edb_top_inst/n740 , \edb_top_inst/n738 , 
        \edb_top_inst/n736 , \edb_top_inst/n734 , \edb_top_inst/n733 , 
        \edb_top_inst/edb_user_dr[65] , \edb_top_inst/edb_user_dr[66] , 
        \edb_top_inst/edb_user_dr[67] , \edb_top_inst/edb_user_dr[68] , 
        \edb_top_inst/edb_user_dr[69] , \edb_top_inst/edb_user_dr[70] , 
        \edb_top_inst/edb_user_dr[71] , \edb_top_inst/edb_user_dr[72] , 
        \edb_top_inst/edb_user_dr[73] , \edb_top_inst/edb_user_dr[74] , 
        \edb_top_inst/edb_user_dr[75] , \edb_top_inst/edb_user_dr[76] , 
        \edb_top_inst/debug_hub_inst/n266 , \edb_top_inst/debug_hub_inst/n95 , 
        \edb_top_inst/edb_user_dr[81] , \edb_top_inst/n714 , \edb_top_inst/n716 , 
        \edb_top_inst/n718 , \edb_top_inst/n720 , \edb_top_inst/n722 , 
        \edb_top_inst/n724 , \edb_top_inst/n726 , \edb_top_inst/n728 , 
        \edb_top_inst/n730 , \edb_top_inst/n732 , \edb_top_inst/n735 , 
        \edb_top_inst/n737 , \edb_top_inst/n739 , \edb_top_inst/n741 , 
        \edb_top_inst/n743 , \edb_top_inst/n745 , \edb_top_inst/n747 , 
        \edb_top_inst/n749 , \edb_top_inst/n751 , \edb_top_inst/n753 , 
        \edb_top_inst/n841 , \edb_top_inst/n843 , \edb_top_inst/n845 , 
        \edb_top_inst/n847 , \edb_top_inst/n849 , \edb_top_inst/n851 , 
        \edb_top_inst/n853 , \edb_top_inst/n855 , \edb_top_inst/n857 , 
        \edb_top_inst/n1009 , \edb_top_inst/n1012 , \edb_top_inst/n1014 , 
        \edb_top_inst/n1016 , \edb_top_inst/n1018 , \edb_top_inst/n1020 , 
        \edb_top_inst/n1022 , \edb_top_inst/n1024 , \edb_top_inst/n1026 , 
        \edb_top_inst/n1029 , \edb_top_inst/n1031 , \edb_top_inst/n1033 , 
        \edb_top_inst/n1035 , \edb_top_inst/n1037 , \edb_top_inst/n1039 , 
        \edb_top_inst/n1041 , \edb_top_inst/n1043 , \edb_top_inst/n1045 , 
        \edb_top_inst/n1048 , \edb_top_inst/n1050 , \edb_top_inst/n1052 , 
        \edb_top_inst/n1065 , \edb_top_inst/n1067 , \edb_top_inst/n1069 , 
        \edb_top_inst/n1071 , \edb_top_inst/n1073 , \edb_top_inst/n1075 , 
        \edb_top_inst/n1077 , \edb_top_inst/n1079 , \edb_top_inst/n1081 , 
        \edb_top_inst/n1083 , \edb_top_inst/n1085 , \edb_top_inst/n1087 , 
        \edb_top_inst/n1089 , \edb_top_inst/n1091 , \edb_top_inst/n1093 , 
        \edb_top_inst/n1095 , \edb_top_inst/n1097 , \edb_top_inst/n1099 , 
        \edb_top_inst/n1101 , \edb_top_inst/n1103 , \edb_top_inst/n1105 , 
        \edb_top_inst/n1107 , \edb_top_inst/n1109 , \edb_top_inst/n1111 , 
        \edb_top_inst/n1113 , \edb_top_inst/n1126 , \edb_top_inst/n1128 , 
        \edb_top_inst/n1130 , \edb_top_inst/n1132 , \edb_top_inst/n1134 , 
        \edb_top_inst/n1136 , \edb_top_inst/n1138 , \edb_top_inst/n1143 , 
        \edb_top_inst/n1145 , \edb_top_inst/n1147 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] , 
        \edb_top_inst/n2758 , \edb_top_inst/n67 , \edb_top_inst/n1112 , 
        \edb_top_inst/n1110 , \edb_top_inst/n1108 , \edb_top_inst/n1106 , 
        \edb_top_inst/n1104 , \edb_top_inst/n1102 , \edb_top_inst/n1100 , 
        \edb_top_inst/n1098 , \edb_top_inst/n1096 , \edb_top_inst/n1094 , 
        \edb_top_inst/n1092 , \edb_top_inst/n1090 , \edb_top_inst/n1088 , 
        \edb_top_inst/n1086 , \edb_top_inst/n1084 , \edb_top_inst/n1082 , 
        \edb_top_inst/n1146 , \edb_top_inst/n1080 , \edb_top_inst/n1144 , 
        \edb_top_inst/n1078 , \edb_top_inst/n1142 , \edb_top_inst/n1076 , 
        \edb_top_inst/n1137 , \edb_top_inst/n1074 , \edb_top_inst/n1135 , 
        \edb_top_inst/n1072 , \edb_top_inst/n1133 , \edb_top_inst/n1070 , 
        \edb_top_inst/n1131 , \edb_top_inst/n1068 , \edb_top_inst/n1129 , 
        \edb_top_inst/n1066 , \edb_top_inst/n1127 , \edb_top_inst/n1064 , 
        \edb_top_inst/n1125 , \edb_top_inst/n1062 , \edb_top_inst/n1123 , 
        \edb_top_inst/n69 , \edb_top_inst/n1051 , \edb_top_inst/n1049 , 
        \edb_top_inst/n1047 , \edb_top_inst/n1046 , \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 , 
        \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 , n8022, n8093, 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5_q , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4_q , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3_q , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2_q , 
        \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1_q , \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0_q , 
        n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, 
        n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, 
        n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, 
        n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, 
        n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, 
        n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, 
        n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, 
        n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, 
        n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, 
        n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, 
        n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, 
        n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, 
        n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, 
        n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, 
        n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, 
        n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, 
        n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, 
        n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, 
        n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8330, 
        n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, 
        n8339, n8340, n8346, n8347, n8348, n8349, n8350, n8351, 
        n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, 
        n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, 
        n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, 
        n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
        n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, 
        n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, 
        n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, 
        n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, 
        n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
        n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, 
        n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, 
        n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, 
        n8448, n8449, n8450, n8451;
    
    assign MipiDphyRx1_RESET_N = MipiDphyRx1_RST0_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[2] = MipiDphyRx1_STOPSTATE_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_REQUEST_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TURN_REQUEST = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_FORCE_RX_MODE = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_TRIGGER_ESC[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[7] = MipiDphyRx1_RX_CLK_ACTIVE_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[10] = MipiDphyRx1_RX_ACTIVE_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[24] = MipiDphyRx1_RX_VALID_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[25] = MipiDphyRx1_RX_VALID_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[0] = MipiDphyRx1_RX_SYNC_HS_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[3] = MipiDphyRx1_RX_SKEW_CAL_HS_LAN1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[4] = MipiDphyRx1_RX_DATA_HS_LAN0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_LPDT_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_DATA_ESC[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_VALID_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_READY_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_ULPS_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign MipiDphyRx1_TX_ULPS_EXIT = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[17] = MipiDphyRx1_WORD_CLKOUT_HS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign oTestPort[1] = MipiDphyRx1_RX_CLK_ESC_LAN0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign MipiDphyRx1_TX_CLK_ESC = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign pll_inst1_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[23] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[22] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[21] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[20] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[19] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[18] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[16] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[15] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[14] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[13] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[12] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[11] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[9] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[8] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign oTestPort[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign jtag_inst1_TDO = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign pll_inst2_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_CELL_NAME=VCC */ ;
    assign oTestPort[5] = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 LUT__11265 (.I0(\la0_probe6[0] ), .I1(oTestPort[24]), .O(\MCsiRxController/n281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11265.LUTMASK = 16'h4444;
    EFX_FF \la0_probe10~FF  (.D(oTestPort[10]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(la0_probe10)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(289)
    defparam \la0_probe10~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe10~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe10~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe10~FF .D_POLARITY = 1'b1;
    defparam \la0_probe10~FF .SR_SYNC = 1'b0;
    defparam \la0_probe10~FF .SR_VALUE = 1'b0;
    defparam \la0_probe10~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe2~FF  (.D(MipiDphyRx1_STOPSTATE_LAN0), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(la0_probe2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(286)
    defparam \la0_probe2~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe2~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe2~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe2~FF .D_POLARITY = 1'b1;
    defparam \la0_probe2~FF .SR_SYNC = 1'b0;
    defparam \la0_probe2~FF .SR_VALUE = 1'b0;
    defparam \la0_probe2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MipiDphyRx1_RESET_N~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iSCLK), 
           .SR(iPushSw[0]), .Q(MipiDphyRx1_RST0_N)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(149)
    defparam \MipiDphyRx1_RESET_N~FF .CLK_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RESET_N~FF .CE_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RESET_N~FF .SR_POLARITY = 1'b0;
    defparam \MipiDphyRx1_RESET_N~FF .D_POLARITY = 1'b1;
    defparam \MipiDphyRx1_RESET_N~FF .SR_SYNC = 1'b0;
    defparam \MipiDphyRx1_RESET_N~FF .SR_VALUE = 1'b0;
    defparam \MipiDphyRx1_RESET_N~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rFRST~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iFCLK), .SR(iPushSw[0]), 
           .Q(rFRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(167)
    defparam \rFRST~FF .CLK_POLARITY = 1'b1;
    defparam \rFRST~FF .CE_POLARITY = 1'b1;
    defparam \rFRST~FF .SR_POLARITY = 1'b0;
    defparam \rFRST~FF .D_POLARITY = 1'b0;
    defparam \rFRST~FF .SR_SYNC = 1'b0;
    defparam \rFRST~FF .SR_VALUE = 1'b1;
    defparam \rFRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rBRST~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iBCLK), .SR(iPushSw[0]), 
           .Q(rBRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(178)
    defparam \rBRST~FF .CLK_POLARITY = 1'b1;
    defparam \rBRST~FF .CE_POLARITY = 1'b1;
    defparam \rBRST~FF .SR_POLARITY = 1'b0;
    defparam \rBRST~FF .D_POLARITY = 1'b0;
    defparam \rBRST~FF .SR_SYNC = 1'b0;
    defparam \rBRST~FF .SR_VALUE = 1'b1;
    defparam \rBRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rVRST~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iVCLK), .SR(iPushSw[0]), 
           .Q(rVRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(189)
    defparam \rVRST~FF .CLK_POLARITY = 1'b1;
    defparam \rVRST~FF .CE_POLARITY = 1'b1;
    defparam \rVRST~FF .SR_POLARITY = 1'b0;
    defparam \rVRST~FF .D_POLARITY = 1'b0;
    defparam \rVRST~FF .SR_SYNC = 1'b0;
    defparam \rVRST~FF .SR_VALUE = 1'b1;
    defparam \rVRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rnVRST~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iVCLK), .SR(iPushSw[0]), 
           .Q(rnVRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(193)
    defparam \rnVRST~FF .CLK_POLARITY = 1'b1;
    defparam \rnVRST~FF .CE_POLARITY = 1'b1;
    defparam \rnVRST~FF .SR_POLARITY = 1'b0;
    defparam \rnVRST~FF .D_POLARITY = 1'b1;
    defparam \rnVRST~FF .SR_SYNC = 1'b0;
    defparam \rnVRST~FF .SR_VALUE = 1'b0;
    defparam \rnVRST~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[2]~FF  (.D(1'b1), .CE(wCdcFifoFull), .CLK(iSCLK), .SR(rSRST), 
           .Q(oLed[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(403)
    defparam \oLed[2]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[2]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[2]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[2]~FF .D_POLARITY = 1'b1;
    defparam \oLed[2]~FF .SR_SYNC = 1'b1;
    defparam \oLed[2]~FF .SR_VALUE = 1'b0;
    defparam \oLed[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe11~FF  (.D(oTestPort[24]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(la0_probe11)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(283)
    defparam \la0_probe11~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe11~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe11~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe11~FF .D_POLARITY = 1'b1;
    defparam \la0_probe11~FF .SR_SYNC = 1'b0;
    defparam \la0_probe11~FF .SR_VALUE = 1'b0;
    defparam \la0_probe11~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[0]~FF  (.D(\MCsiRxController/n281 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[0]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[0]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(280)
    defparam \la0_probe9[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/n631 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/n633 ), 
           .Q(\MCsiRxController/MCsi2Decoder/rHsSt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(213)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe3[0]~FF  (.D(oTestPort[0]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe3[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe3[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe3[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe3[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe3[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe3[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe3[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe3[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF  (.D(\MCsiRxController/MCsi2Decoder/n7 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rSRST_2~FF  (.D(oLed[5]), .CE(1'b1), .CLK(iSCLK), .SR(iPushSw[0]), 
           .Q(rSRST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MTopTi180MIPI25GRxHDMIV101.v(145)
    defparam \rSRST_2~FF .CLK_POLARITY = 1'b1;
    defparam \rSRST_2~FF .CE_POLARITY = 1'b1;
    defparam \rSRST_2~FF .SR_POLARITY = 1'b0;
    defparam \rSRST_2~FF .D_POLARITY = 1'b0;
    defparam \rSRST_2~FF .SR_SYNC = 1'b0;
    defparam \rSRST_2~FF .SR_VALUE = 1'b1;
    defparam \rSRST_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe4~FF  (.D(MipiDphyRx1_RX_SKEW_CAL_HS_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(la0_probe4)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(292)
    defparam \la0_probe4~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe4~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe4~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe4~FF .D_POLARITY = 1'b1;
    defparam \la0_probe4~FF .SR_SYNC = 1'b0;
    defparam \la0_probe4~FF .SR_VALUE = 1'b0;
    defparam \la0_probe4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe5~FF  (.D(MipiDphyRx1_ERR_SOT_HS_LAN0), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(la0_probe5)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(295)
    defparam \la0_probe5~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe5~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe5~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe5~FF .D_POLARITY = 1'b1;
    defparam \la0_probe5~FF .SR_SYNC = 1'b0;
    defparam \la0_probe5~FF .SR_VALUE = 1'b0;
    defparam \la0_probe5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe7~FF  (.D(MipiDphyRx1_RX_ERR_SYNC_ESC), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(la0_probe7)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(298)
    defparam \la0_probe7~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe7~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe7~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe7~FF .D_POLARITY = 1'b1;
    defparam \la0_probe7~FF .SR_SYNC = 1'b0;
    defparam \la0_probe7~FF .SR_VALUE = 1'b0;
    defparam \la0_probe7~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe0~FF  (.D(la0_probe0), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(la0_probe0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(268)
    defparam \la0_probe0~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe0~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe0~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe0~FF .D_POLARITY = 1'b0;
    defparam \la0_probe0~FF .SR_SYNC = 1'b0;
    defparam \la0_probe0~FF .SR_VALUE = 1'b0;
    defparam \la0_probe0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(115)
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiRvd[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wCddFifoFull~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qFullAllmost ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(wCddFifoFull)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(105)
    defparam \wCddFifoFull~FF .CLK_POLARITY = 1'b1;
    defparam \wCddFifoFull~FF .CE_POLARITY = 1'b1;
    defparam \wCddFifoFull~FF .SR_POLARITY = 1'b0;
    defparam \wCddFifoFull~FF .D_POLARITY = 1'b1;
    defparam \wCddFifoFull~FF .SR_SYNC = 1'b0;
    defparam \wCddFifoFull~FF .SR_VALUE = 1'b0;
    defparam \wCddFifoFull~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsValid~FF  (.D(\MCsiRxController/MCsi2Decoder/n585 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsValid )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsValid~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/wHsValid~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsValid~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsValid~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/n97 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(rSRST), .Q(\MCsiRxController/MCsi2Decoder/rHsSt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(213)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/n607 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/n633 ), 
           .Q(\MCsiRxController/MCsi2Decoder/rHsSt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(213)
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rHsSt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[7]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[7]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe9[7]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[7]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[7]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[7]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[7]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[7]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[6]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[6]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe9[6]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[6]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[6]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[6]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[6]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[6]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[5]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[5]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe9[5]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[5]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[5]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[5]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[5]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[5]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[4]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[4]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe9[4]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[4]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[4]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[4]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[4]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[4]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[3]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[3]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe9[3]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[3]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[3]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[3]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[3]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[3]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[2]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[2]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe9[2]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[2]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[2]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[2]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[2]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[2]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe9[1]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN1[1]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe9[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe9[1]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe9[1]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe9[1]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe9[1]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe9[1]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe9[1]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe9[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n19 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/wFtiEmp[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(112)
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_VALUE = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/wFtiEmp[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF  (.D(n116), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF  (.D(n3019), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF  (.D(n3017), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF  (.D(n3015), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF  (.D(n3013), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF  (.D(n3011), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF  (.D(n3009), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF  (.D(n3007), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF  (.D(n3006), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n233 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n238 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n243 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n248 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n253 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n258 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n263 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n268 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n273 ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd ), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF  (.D(n119), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF  (.D(n169), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF  (.D(n2983), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF  (.D(n2981), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF  (.D(n2979), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF  (.D(n2977), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF  (.D(n2975), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF  (.D(n2973), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF  (.D(n2972), 
           .CE(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[9] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[10]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[10] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[11]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[11] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[12]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[12] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[13]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[13] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[13]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[14]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[14] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[14]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wHsPixel[15]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[15] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(1'b0), .Q(\MCsiRxController/wHsPixel[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/wHsPixel[15]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/wHsPixel[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[1]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[9] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[10] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[11] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[12] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[13] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[6]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[14] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[7]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[15] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[8]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[0] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_60/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[9]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[1] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_60/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[10]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_60/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[11]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_60/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[11]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[11]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[12]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_60/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[12]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[12]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[13]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_60/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[13]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[13]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[13]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[14]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[6] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_60/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[14]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[14]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[14]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsWordCnt[15]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[7] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_60/n5 ), .CLK(iSCLK), 
           .SR(1'b0), .Q(\wHsWordCnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsWordCnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .CE_POLARITY = 1'b0;
    defparam \wHsWordCnt[15]~FF .SR_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .D_POLARITY = 1'b1;
    defparam \wHsWordCnt[15]~FF .SR_SYNC = 1'b1;
    defparam \wHsWordCnt[15]~FF .SR_VALUE = 1'b0;
    defparam \wHsWordCnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[2]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[2] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsDatatype[2]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[2]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[2]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[2]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[3]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[3] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsDatatype[3]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[3]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[3]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[3]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[4]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[4] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsDatatype[4]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[4]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[4]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[4]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wHsDatatype[5]~FF  (.D(\MCsiRxController/MCsi2Decoder/wFtiRd[5] ), 
           .CE(\MCsiRxController/MCsi2Decoder/equal_63/n5 ), .CLK(iSCLK), 
           .SR(rSRST), .Q(\wHsDatatype[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \wHsDatatype[5]~FF .CLK_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .CE_POLARITY = 1'b0;
    defparam \wHsDatatype[5]~FF .SR_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .D_POLARITY = 1'b1;
    defparam \wHsDatatype[5]~FF .SR_SYNC = 1'b1;
    defparam \wHsDatatype[5]~FF .SR_VALUE = 1'b0;
    defparam \wHsDatatype[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF  (.D(n124), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF  (.D(n3004), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF  (.D(n3002), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF  (.D(n3000), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF  (.D(n2998), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF  (.D(n2996), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF  (.D(n2994), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF  (.D(n2992), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF  (.D(n2990), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF  (.D(n2988), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF  (.D(n2986), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF  (.D(n2985), 
           .CE(\MCsiRxController/MCsi2Decoder/n604 ), .CLK(iSCLK), .SR(\MCsiRxController/MCsi2Decoder/qLineCntRst ), 
           .Q(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(274)
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_SYNC = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[0]~FF  (.D(oTestPort[4]), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe8[0]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[0]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[0]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[0]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[0]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[0]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[1]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[1]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe8[1]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[1]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[1]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[1]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[1]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[1]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[2]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[2]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe8[2]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[2]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[2]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[2]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[2]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[2]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[3]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[3]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe8[3]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[3]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[3]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[3]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[3]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[3]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[4]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[4]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe8[4]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[4]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[4]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[4]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[4]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[4]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[5]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[5]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe8[5]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[5]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[5]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[5]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[5]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[5]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[6]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[6]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe8[6]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[6]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[6]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[6]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[6]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[6]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe8[7]~FF  (.D(MipiDphyRx1_RX_DATA_HS_LAN0[7]), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe8[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(127)
    defparam \la0_probe8[7]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe8[7]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe8[7]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe8[7]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe8[7]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe8[7]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe8[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wCdcFifoFull_2~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(wCdcFifoFull)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(85)
    defparam \wCdcFifoFull_2~FF .CLK_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .CE_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .SR_POLARITY = 1'b0;
    defparam \wCdcFifoFull_2~FF .D_POLARITY = 1'b1;
    defparam \wCdcFifoFull_2~FF .SR_SYNC = 1'b0;
    defparam \wCdcFifoFull_2~FF .SR_VALUE = 1'b0;
    defparam \wCdcFifoFull_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wVideoVd~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/qRVD ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(wVideoVd)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(91)
    defparam \wVideoVd~FF .CLK_POLARITY = 1'b1;
    defparam \wVideoVd~FF .CE_POLARITY = 1'b1;
    defparam \wVideoVd~FF .SR_POLARITY = 1'b0;
    defparam \wVideoVd~FF .D_POLARITY = 1'b1;
    defparam \wVideoVd~FF .SR_SYNC = 1'b0;
    defparam \wVideoVd~FF .SR_VALUE = 1'b0;
    defparam \wVideoVd~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/wFtiEmp[0]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/wFtiEmp[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(88)
    defparam \MCsiRxController/wFtiEmp[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .D_POLARITY = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_VALUE = 1'b1;
    defparam \MCsiRxController/wFtiEmp[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF  (.D(n189), .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF  (.D(n210), .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), 
           .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF  (.D(n2970), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF  (.D(n2968), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF  (.D(n2966), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF  (.D(n2964), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF  (.D(n2962), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF  (.D(n2961), 
           .CE(\MCsiRxController/genblk1[0].mVideoFIFO/qRE ), .CLK(iSCLK), 
           .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(64)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rRA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(67)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n436 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n441 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n446 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n451 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n456 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n461 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n466 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF  (.D(\MCsiRxController/genblk1[0].mVideoFIFO/n471 ), 
           .CE(\MCsiRxController/wHsValid ), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), 
           .Q(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(60)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[1]~FF  (.D(\MCsiRxController/n280 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[1]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[1]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[1]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[1]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[1]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[1]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[2]~FF  (.D(\MCsiRxController/n279 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[2]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[2]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[2]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[2]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[2]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[2]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[3]~FF  (.D(\MCsiRxController/n278 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[3]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[3]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[3]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[3]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[3]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[3]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[4]~FF  (.D(\MCsiRxController/n277 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[4]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[4]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[4]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[4]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[4]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[4]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[5]~FF  (.D(\MCsiRxController/n276 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[5]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[5]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[5]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[5]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[5]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[5]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[6]~FF  (.D(\MCsiRxController/n275 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[6]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[6]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[6]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[6]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[6]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[6]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[7]~FF  (.D(\MCsiRxController/n274 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[7]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[7]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[7]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[7]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[7]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[7]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[8]~FF  (.D(\MCsiRxController/n273 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[8]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[8]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[8]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[8]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[8]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[8]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[9]~FF  (.D(\MCsiRxController/n272 ), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[9]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[9]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[9]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[9]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[9]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[9]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[10]~FF  (.D(\MCsiRxController/n271 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[10]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[10]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[10]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[10]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[10]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[10]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[11]~FF  (.D(\MCsiRxController/n270 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[11]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[11]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[11]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[11]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[11]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[11]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[12]~FF  (.D(\MCsiRxController/n269 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[12]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[12]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[12]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[12]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[12]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[12]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[13]~FF  (.D(\MCsiRxController/n268 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[13]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[13]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[13]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[13]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[13]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[13]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[14]~FF  (.D(\MCsiRxController/n267 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[14]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[14]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[14]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[14]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[14]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[14]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe6[15]~FF  (.D(\MCsiRxController/n266 ), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe6[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(302)
    defparam \la0_probe6[15]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe6[15]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe6[15]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe6[15]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe6[15]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe6[15]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe6[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \la0_probe3[1]~FF  (.D(MipiDphyRx1_RX_SYNC_HS_LAN1), .CE(1'b1), 
           .CLK(oTestPort[17]), .SR(MipiDphyRx1_RST0_N), .Q(\la0_probe3[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(274)
    defparam \la0_probe3[1]~FF .CLK_POLARITY = 1'b1;
    defparam \la0_probe3[1]~FF .CE_POLARITY = 1'b1;
    defparam \la0_probe3[1]~FF .SR_POLARITY = 1'b0;
    defparam \la0_probe3[1]~FF .D_POLARITY = 1'b1;
    defparam \la0_probe3[1]~FF .SR_SYNC = 1'b0;
    defparam \la0_probe3[1]~FF .SR_VALUE = 1'b0;
    defparam \la0_probe3[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[0]~FF  (.D(\MVideoPostProcess/rVtgRstCnt[0] ), 
           .CE(\MVideoPostProcess/qVtgRstCntCke ), .CLK(iVCLK), .SR(rVRST), 
           .Q(\MVideoPostProcess/rVtgRstCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[0]~FF  (.D(\MVideoPostProcess/rVtgRstSel ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRST[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstSel_2~FF  (.D(1'b0), .CE(\MVideoPostProcess/equal_18/n21 ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstSel )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRstSel_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF  (.D(\~n1835 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n816 ), 
           .CE(\~ceg_net512 ), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_m_en_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n833 ), 
           .CE(\~ceg_net512 ), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_last_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_last_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n268 ), 
           .CE(ceg_net995), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n277 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF  (.D(ceg_net43), 
           .CE(ceg_net1327), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1243 ), .CLK(iBCLK), 
           .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1243 ), .CLK(iBCLK), 
           .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_3P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 ), 
           .CE(ceg_net1087), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511SdaOe~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 ), 
           .CE(ceg_net1335), .CLK(iBCLK), .SR(rBRST), .Q(oAdv7511SdaOe)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \oAdv7511SdaOe~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .CE_POLARITY = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511SdaOe~FF .SR_SYNC = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511SdaOe~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511SclOe~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 ), 
           .CE(ceg_net566), .CLK(iBCLK), .SR(rBRST), .Q(oAdv7511SclOe)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \oAdv7511SclOe~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .CE_POLARITY = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511SclOe~FF .SR_SYNC = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511SclOe~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 ), 
           .CE(ceg_net1361), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/w_ack~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/w_ack )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/w_ack~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 ), 
           .CE(ceg_net616), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 ), 
           .CE(1'b1), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 ), 
           .CE(ceg_net1087), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 ), 
           .CE(ceg_net1087), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 ), 
           .CE(ceg_net1400), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 ), 
           .CE(ceg_net1463), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 ), 
           .CE(ceg_net1471), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 ), 
           .CE(ceg_net1480), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 ), 
           .CE(ceg_net1488), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\i2c_phy.v(677)
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n8455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4659)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(1'b1), .CI(1'b0), .CO(n8454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4673)
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4  (.I0(n8093), 
            .I1(1'b1), .CI(1'b0), .CO(n8453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__MVideoPostProcess/mVideoTimingGen/add_6/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0_q ), 
            .I1(1'b1), .CI(1'b0), .CO(n8452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n251 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n250 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n249 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n248 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n247 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n246 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n245 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n244 ), 
           .CE(ceg_net939), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_addr_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n700 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n705 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n710 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n715 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n720 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n725 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n730 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n735 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n740 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n745 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n750 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n755 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n760 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n765 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n770 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1107 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n780 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n785 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n790 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n795 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n800 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n805 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n810 ), 
           .CE(\MVideoPostProcess/inst_adv7511_config/n1224 ), .CLK(iBCLK), 
           .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n276 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n275 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n274 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n273 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n272 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n271 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/n270 ), 
           .CE(ceg_net479), .CLK(iBCLK), .SR(1'b0), .Q(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF  (.D(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
           .CE(ceg_net1327), .CLK(iBCLK), .SR(rBRST), .Q(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\sample\adv7511_config.v(279)
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n131 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/qVde ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rVde[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511Hs~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rHSync[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511Hs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \oAdv7511Hs~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511Hs~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511Hs~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511Hs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n130 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n129 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF  (.D(n2917), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF  (.D(n2915), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n126 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n125 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF  (.D(n2909), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF  (.D(n2907), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF  (.D(n2905), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/n121 ), 
           .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), .CLK(iVCLK), 
           .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF  (.D(n2902), .CE(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), .Q(\MVideoPostProcess/mVideoTimingGen/rVpos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .CE_POLARITY = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVpos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511Vs~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVSync[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511Vs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \oAdv7511Vs~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511Vs~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511Vs~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511Vs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVde[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rVde[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF  (.D(\MVideoPostProcess/wVgaGenFDe ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/rVde[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rVde[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oAdv7511De~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVde[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(oAdv7511De)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \oAdv7511De~FF .CLK_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .CE_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .SR_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .D_POLARITY = 1'b1;
    defparam \oAdv7511De~FF .SR_SYNC = 1'b1;
    defparam \oAdv7511De~FF .SR_VALUE = 1'b0;
    defparam \oAdv7511De~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/wVgaGenFDe_2~FF  (.D(\MVideoPostProcess/mVideoTimingGen/rVde[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/wVgaGenFDe )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(120)
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/wVgaGenFDe_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF  (.D(n436), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF  (.D(n2938), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF  (.D(n2936), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF  (.D(n2934), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF  (.D(n2932), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF  (.D(n2930), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF  (.D(n2928), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF  (.D(n2926), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF  (.D(n2924), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF  (.D(n2922), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF  (.D(n2921), .CE(1'b1), 
           .CLK(iVCLK), .SR(\MVideoPostProcess/mVideoTimingGen/n267 ), .Q(\MVideoPostProcess/mVideoTimingGen/rHpos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/mVideoTimingGen/rHpos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \wVideofull~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost ), 
           .CE(1'b1), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(wVideofull)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(105)
    defparam \wVideofull~FF .CLK_POLARITY = 1'b1;
    defparam \wVideofull~FF .CE_POLARITY = 1'b1;
    defparam \wVideofull~FF .SR_POLARITY = 1'b0;
    defparam \wVideofull~FF .D_POLARITY = 1'b1;
    defparam \wVideofull~FF .SR_SYNC = 1'b0;
    defparam \wVideofull~FF .SR_VALUE = 1'b0;
    defparam \wVideofull~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n492), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n2900), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n2898), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n2896), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n2894), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n2892), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n2890), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n2888), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n2886), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n2885), 
           .CE(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n433 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n438 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n443 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n448 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n453 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n458 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n463 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n468 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n473 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF  (.D(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n532), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n555), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n2883), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n2881), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n2879), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n2877), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n2875), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n2873), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n2871), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n2870), 
           .CE(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n573), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n596), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n2868), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n2866), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n2864), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n2862), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n2860), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n2858), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n2856), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n2855), 
           .CE(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] ), 
           .CE(wVideoVd), .CLK(iSCLK), .SR(MipiDphyRx1_RST0_N), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(64)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .D_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF  (.D(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(81)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF  (.D(n614), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF  (.D(n637), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF  (.D(n2853), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF  (.D(n2851), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF  (.D(n2849), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF  (.D(n2847), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF  (.D(n2845), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF  (.D(n2843), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF  (.D(n2841), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF  (.D(n2840), 
           .CE(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE ), .CLK(iVCLK), 
           .SR(rnVRST), .Q(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(85)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[1]~FF  (.D(n295), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[2]~FF  (.D(n331), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[3]~FF  (.D(n2959), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[4]~FF  (.D(n2957), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[5]~FF  (.D(n2955), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[6]~FF  (.D(n2953), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[7]~FF  (.D(n2951), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[8]~FF  (.D(n2949), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[9]~FF  (.D(n2947), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRstCnt[10]~FF  (.D(n2946), .CE(\MVideoPostProcess/qVtgRstCntCke ), 
           .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRstCnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_VALUE = 1'b0;
    defparam \MVideoPostProcess/rVtgRstCnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[1]~FF  (.D(\MVideoPostProcess/rVtgRST[0] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRST[1]~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/rVtgRST[2]_2~FF  (.D(\MVideoPostProcess/rVtgRST[1] ), 
           .CE(1'b1), .CLK(iVCLK), .SR(rVRST), .Q(\MVideoPostProcess/rVtgRST[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(189)
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/rVtgRST[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[0]~FF  (.D(oLed[0]), .CE(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), 
           .CLK(iFCLK), .SR(rFRST), .Q(oLed[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(71)
    defparam \oLed[0]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[0]~FF .CE_POLARITY = 1'b0;
    defparam \oLed[0]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[0]~FF .D_POLARITY = 1'b0;
    defparam \oLed[0]~FF .SR_SYNC = 1'b1;
    defparam \oLed[0]~FF .SR_VALUE = 1'b0;
    defparam \oLed[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF  (.D(wVideoVd), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5  (.D(n8022), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5 .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5 .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5 .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5 .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5 .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5 .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF  (.D(n2838), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF  (.D(n2836), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF  (.D(n2834), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF  (.D(n2832), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF  (.D(n2830), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF  (.D(n2828), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF  (.D(n2826), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF  (.D(n2824), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF  (.D(n2823), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[0].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[0].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[1].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[1].mPulseGenerator/equal_12/n3 ), .Q(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[1]~FF  (.D(oLed[1]), .CE(\genblk1.genblk1[1].mPulseGenerator/equal_12/n3 ), 
           .CLK(iFCLK), .SR(rFRST), .Q(oLed[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(71)
    defparam \oLed[1]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[1]~FF .CE_POLARITY = 1'b0;
    defparam \oLed[1]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[1]~FF .D_POLARITY = 1'b0;
    defparam \oLed[1]~FF .SR_SYNC = 1'b1;
    defparam \oLed[1]~FF .SR_VALUE = 1'b0;
    defparam \oLed[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF  (.D(wCddFifoFull), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[1].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF  (.D(\genblk1.genblk1[1].mPulseGenerator/n50 ), 
           .CE(\genblk1.genblk1[1].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[1].mPulseGenerator/equal_12/n3 ), .Q(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[1].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[1].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[1].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[1].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[1].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[3]~FF  (.D(oLed[3]), .CE(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), 
           .CLK(iFCLK), .SR(rFRST), .Q(oLed[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(71)
    defparam \oLed[3]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[3]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[3]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[3]~FF .D_POLARITY = 1'b0;
    defparam \oLed[3]~FF .SR_SYNC = 1'b1;
    defparam \oLed[3]~FF .SR_VALUE = 1'b0;
    defparam \oLed[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF  (.D(wCdcFifoFull), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/n50 ), 
           .CE(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[3].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[3].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[3].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] ), 
           .CE(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .D_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \oLed[4]~FF  (.D(oLed[4]), .CE(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), 
           .CLK(iFCLK), .SR(rFRST), .Q(oLed[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(71)
    defparam \oLed[4]~FF .CLK_POLARITY = 1'b1;
    defparam \oLed[4]~FF .CE_POLARITY = 1'b1;
    defparam \oLed[4]~FF .SR_POLARITY = 1'b1;
    defparam \oLed[4]~FF .D_POLARITY = 1'b0;
    defparam \oLed[4]~FF .SR_SYNC = 1'b1;
    defparam \oLed[4]~FF .SR_VALUE = 1'b0;
    defparam \oLed[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF  (.D(wVideofull), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/n50 ), 
           .CE(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .Q(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rTmpCount[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rSft[0] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF  (.D(\genblk1.genblk1[4].mPulseGenerator/rSft[1] ), 
           .CE(1'b1), .CLK(iFCLK), .SR(rFRST), .Q(\genblk1.genblk1[4].mPulseGenerator/rSft[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(36)
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .CE_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[4].mPulseGenerator/rSft[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(69)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_2_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF  (.D(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_rst_0 ), 
           .CE(1'b1), .CLK(iVCLK), .SR(\MVideoPostProcess/rVtgRST[2] ), 
           .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(97)
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .CE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .D_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_SYNC = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_VALUE = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_1_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n1340 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1341 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1342 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n1965 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3683)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[0] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n2189 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[0] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2466 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state[0] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3794)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_soft_reset_in ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4104)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_soft_reset_in ), 
           .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4104)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(la0_probe0), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(la0_probe1), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF  (.D(la0_probe2), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF  (.D(\la0_probe3[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5294 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5492 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF  (.D(la0_probe4), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF  (.D(la0_probe5), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6947 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF  (.D(\la0_probe6[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF  (.D(la0_probe7), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n8741 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF  (.D(\la0_probe8[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF  (.D(\la0_probe9[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10527 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF  (.D(la0_probe10), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n11368 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF  (.D(la0_probe11), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n12201 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1396 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3656)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1913 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3668)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[1] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[2] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[3] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[4] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[5] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[6] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[7] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[8] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[9] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[10] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[11] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[12] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[13] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[14] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[15] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[16] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[17] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[18] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[19] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[20] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[21] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[22] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[23] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[24] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[25]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[25] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[26]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[26] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/address_counter[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3702)
    defparam \edb_top_inst/la0/address_counter[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/opcode[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n2188 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n2187 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n2186 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n2185 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n2184 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/bit_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[1] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[2] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[3] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[4] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[5] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[6] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[7] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[8] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[9] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[10] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[11] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[12] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[13] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[14] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[15] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/word_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3739)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2465 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2464 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2463 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2462 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2461 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2460 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2459 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2458 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2457 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2456 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2455 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2454 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2453 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2452 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2451 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2450 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2449 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2448 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2447 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2446 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2445 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2444 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2443 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2442 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2441 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2440 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2439 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2438 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2437 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2436 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2435 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2434 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2433 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2432 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2431 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2430 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2429 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2428 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2427 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2426 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2425 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2424 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2423 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2422 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2421 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2420 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2419 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2418 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2417 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2416 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2415 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2414 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2413 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2412 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2411 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2410 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2409 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2408 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2407 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2406 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2405 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2404 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2403 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3752)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state[1] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3794)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state[2] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3794)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state[3] ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/module_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3794)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n150 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n149 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n148 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n147 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n146 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n145 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n144 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n143 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n142 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n141 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n140 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n139 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n138 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n137 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n136 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n135 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n134 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n133 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n132 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n131 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n130 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n129 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n128 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n127 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n126 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n125 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n124 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n123 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n122 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n121 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n120 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n119 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(284)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2766 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2766 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n2766 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5522)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3599 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3599 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3599 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4432 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4432 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4432 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF  (.D(\la0_probe3[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5279 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5279 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5279 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5294 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5492 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n10 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n3 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n9 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6114 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6114 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6114 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6947 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6947 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF  (.D(\la0_probe6[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF  (.D(\la0_probe6[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF  (.D(\la0_probe6[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF  (.D(\la0_probe6[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF  (.D(\la0_probe6[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF  (.D(\la0_probe6[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF  (.D(\la0_probe6[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF  (.D(\la0_probe6[8] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF  (.D(\la0_probe6[9] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF  (.D(\la0_probe6[10] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF  (.D(\la0_probe6[11] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF  (.D(\la0_probe6[12] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF  (.D(\la0_probe6[13] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF  (.D(\la0_probe6[14] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF  (.D(\la0_probe6[15] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7892 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7892 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7892 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n7907 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n8105 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n72 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n73 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n31 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n82 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n71 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n32 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n31 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n30 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n29 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n28 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n27 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n26 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n25 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n24 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n8741 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n8741 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF  (.D(\la0_probe8[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF  (.D(\la0_probe8[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF  (.D(\la0_probe8[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF  (.D(\la0_probe8[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF  (.D(\la0_probe8[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF  (.D(\la0_probe8[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF  (.D(\la0_probe8[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n9630 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9630 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9630 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n9645 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n9843 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF  (.D(\la0_probe9[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF  (.D(\la0_probe9[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF  (.D(\la0_probe9[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF  (.D(\la0_probe9[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF  (.D(\la0_probe9[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF  (.D(\la0_probe9[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF  (.D(\la0_probe9[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4131)
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n21 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n20 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10527 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10527 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n10542 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n10740 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n21 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5634)
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n11368 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n11368 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n12201 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n12201 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5583)
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n89 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5764)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[40]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[41]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4428)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[23] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[40]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[40] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[41]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[41] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4440)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5250)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5050)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5050)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5050)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5271)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5286)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5286)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5286)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5296)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5309)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5309)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5309)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5433)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1300 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/n17781 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5250)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5250)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5250)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5050)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n382 ), 
           .CE(\edb_top_inst/ceg_net348 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5321)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF  (.D(\edb_top_inst/la0/address_counter[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF  (.D(\edb_top_inst/la0/address_counter[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n382 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5331)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[1] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[2] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[5] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[6] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[7] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[8] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[9] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[10] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[11] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[12] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[13]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[13] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[14]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[14] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[15]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[16]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[17]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[18]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[19]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[20]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[21]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[22]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[23]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[24]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[25]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[26]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[27]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[27] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[28]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[28] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[29]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[29] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[30]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[30] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[31]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[31] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[32]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[32] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[33]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[33] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[34]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[34] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[35]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[35] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[36]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[36] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[37]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[37] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[38]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[38] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[39]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[39] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[40]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[40] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[41]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[41] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[42]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[42] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1315 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5340)
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(5433)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/n2053 ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/n73 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/n1044 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/n1042 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/n1040 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/n1038 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/n1036 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/n1034 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/n1032 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/n1030 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF  (.D(\edb_top_inst/n1028 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF  (.D(\edb_top_inst/n1027 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/n693 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/n1025 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/n1023 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/n1021 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/n1019 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/n1017 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/n1015 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/n1013 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/n1011 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF  (.D(\edb_top_inst/n1008 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF  (.D(\edb_top_inst/n1005 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n2053 ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/n695 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/n856 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/n854 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/n852 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/n850 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/n848 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/n846 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/n844 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/n842 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF  (.D(\edb_top_inst/n840 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF  (.D(\edb_top_inst/n838 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(oTestPort[17]), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/n710 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/n731 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/n729 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/n727 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/n725 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/n723 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/n721 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/n719 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/n717 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/n715 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[11]~FF  (.D(\edb_top_inst/n713 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[12]~FF  (.D(\edb_top_inst/n712 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4680)
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[23] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[40] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[41] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4749)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] ), 
           .CE(1'b1), .CLK(oTestPort[17]), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4571)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/n711 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/n752 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/n750 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/n748 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/n746 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/n744 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/n742 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/n740 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/n738 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF  (.D(\edb_top_inst/n736 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF  (.D(\edb_top_inst/n734 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF  (.D(\edb_top_inst/n733 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(oTestPort[17]), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4666)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/internal_register_select[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3597)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1312 ), .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3646)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(355)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]_2~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(355)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(355)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(355)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]_2~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]_2~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]_2~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]_2~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]_2~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]_2~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]_2~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]_2~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]_2~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]_2~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]_2~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]_2~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]_2~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]_2~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]_2~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]_2~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]_2~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]_2~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]_2~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]_2~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]_2~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]_2~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]_2~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]_2~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]_2~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]_2~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]_2~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]_2~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]_2~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]_2~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]_2~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]_2~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]_2~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]_2~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]_2~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]_2~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]_2~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]_2~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]_2~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]_2~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]_2~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]_2~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]_2~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]_2~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]_2~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]_2~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]_2~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]_2~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]_2~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]_2~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]_2~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]_2~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]_2~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]_2~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]_2~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]_2~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]_2~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]_2~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]_2~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]_2~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]_2~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]_2~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]_2~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]_2~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]_2~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]_2~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]_2~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]_2~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]_2~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]_2~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]_2~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]_2~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]_2~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]_2~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]_2~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]_2~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]_2~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]_2~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]_2~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]_2~FF  (.D(\edb_top_inst/edb_user_dr[81] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(jtag_inst2_TCK), 
           .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]_2~FF  (.D(jtag_inst2_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(jtag_inst2_TCK), .SR(jtag_inst2_RESET), .Q(\edb_top_inst/edb_user_dr[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(348)
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .CI(1'b0), .O(n116), .CO(n117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i2  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] ), 
            .CI(1'b0), .O(n119), .CO(n120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i2  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), .CI(1'b0), 
            .O(n124), .CO(n125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i3  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(1'b0), .CI(n120), .O(n169), .CO(n170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), .CI(1'b0), 
            .O(n189), .CO(n190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n190), .O(n210), .CO(n211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i2  (.I0(\MVideoPostProcess/rVtgRstCnt[1] ), 
            .I1(\MVideoPostProcess/rVtgRstCnt[0] ), .CI(1'b0), .O(n295), 
            .CO(n296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i3  (.I0(\MVideoPostProcess/rVtgRstCnt[2] ), 
            .I1(1'b0), .CI(n296), .O(n331), .CO(n332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i2  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[1] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), .CI(1'b0), 
            .O(n436), .CO(n437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i2  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[1] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), .CI(1'b0), 
            .O(n489), .CO(n490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n492), .CO(n493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n532), .CO(n533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n533), .O(n555), .CO(n556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n573), .CO(n574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n574), .O(n596), .CO(n597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
            .CI(1'b0), .O(n614), .CO(n615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n615), .O(n637), .CO(n638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i2  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3_q ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), .CI(1'b0), 
            .O(n655), .CO(n656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i2 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i3  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4_q ), 
            .I1(1'b0), .CI(n656), .O(n678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i3 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i12  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[11] ), 
            .I1(1'b0), .CI(n2825), .O(n2823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i12 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i11  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[10] ), 
            .I1(1'b0), .CI(n2827), .O(n2824), .CO(n2825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i11 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i10  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[9] ), 
            .I1(1'b0), .CI(n2829), .O(n2826), .CO(n2827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i10 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i9  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8] ), 
            .I1(1'b0), .CI(n2831), .O(n2828), .CO(n2829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i9 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i8  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] ), 
            .I1(1'b0), .CI(n2833), .O(n2830), .CO(n2831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i8 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i7  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[6] ), 
            .I1(1'b0), .CI(n2835), .O(n2832), .CO(n2833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i7 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i6  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5] ), 
            .I1(1'b0), .CI(n2837), .O(n2834), .CO(n2835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i6 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i5  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[4] ), 
            .I1(1'b0), .CI(n2839), .O(n2836), .CO(n2837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i5 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \genblk1.genblk1[0].mPulseGenerator/add_8/i4  (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] ), 
            .I1(1'b0), .CI(n8452), .O(n2838), .CO(n2839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(52)
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n2842), .O(n2840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n2844), .O(n2841), .CO(n2842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n2846), .O(n2843), .CO(n2844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n2848), .O(n2845), .CO(n2846)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n2850), .O(n2847), .CO(n2848)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n2852), .O(n2849), .CO(n2850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n2854), .O(n2851), .CO(n2852)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n638), .O(n2853), .CO(n2854)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n2857), .O(n2855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n2859), .O(n2856), .CO(n2857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n2861), .O(n2858), .CO(n2859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n2863), .O(n2860), .CO(n2861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n2865), .O(n2862), .CO(n2863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n2867), .O(n2864), .CO(n2865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n2869), .O(n2866), .CO(n2867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n597), .O(n2868), .CO(n2869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n2872), .O(n2870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n2874), .O(n2871), .CO(n2872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n2876), .O(n2873), .CO(n2874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n2878), .O(n2875), .CO(n2876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n2880), .O(n2877), .CO(n2878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n2882), .O(n2879), .CO(n2880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n2884), .O(n2881), .CO(n2882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n556), .O(n2883), .CO(n2884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(1'b0), .CI(n2887), .O(n2885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
            .I1(1'b0), .CI(n2889), .O(n2886), .CO(n2887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n2891), .O(n2888), .CO(n2889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n2893), .O(n2890), .CO(n2891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n2895), .O(n2892), .CO(n2893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n2897), .O(n2894), .CO(n2895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n2899), .O(n2896), .CO(n2897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n2901), .O(n2898), .CO(n2899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3  (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .I1(1'b0), .CI(n493), .O(n2900), .CO(n2901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i12  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I1(1'b0), .CI(n2904), .O(n2902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i11  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I1(1'b0), .CI(n2906), .O(n2903), .CO(n2904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i10  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[9] ), 
            .I1(1'b0), .CI(n2908), .O(n2905), .CO(n2906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i9  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[8] ), 
            .I1(1'b0), .CI(n2910), .O(n2907), .CO(n2908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i8  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[7] ), 
            .I1(1'b0), .CI(n2912), .O(n2909), .CO(n2910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i7  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), 
            .I1(1'b0), .CI(n2914), .O(n2911), .CO(n2912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i6  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), 
            .I1(1'b0), .CI(n2916), .O(n2913), .CO(n2914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i5  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I1(1'b0), .CI(n2918), .O(n2915), .CO(n2916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i4  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .I1(1'b0), .CI(n2920), .O(n2917), .CO(n2918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_20/i3  (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .I1(1'b0), .CI(n490), .O(n2919), .CO(n2920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(89)
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_20/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i12  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), 
            .I1(1'b0), .CI(n2923), .O(n2921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i12 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i11  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), 
            .I1(1'b0), .CI(n2925), .O(n2922), .CO(n2923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i10  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), 
            .I1(1'b0), .CI(n2927), .O(n2924), .CO(n2925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i9  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), 
            .I1(1'b0), .CI(n2929), .O(n2926), .CO(n2927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i8  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I1(1'b0), .CI(n2931), .O(n2928), .CO(n2929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i7  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I1(1'b0), .CI(n2933), .O(n2930), .CO(n2931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i6  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), 
            .I1(1'b0), .CI(n2935), .O(n2932), .CO(n2933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i5  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), 
            .I1(1'b0), .CI(n2937), .O(n2934), .CO(n2935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i4  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), 
            .I1(1'b0), .CI(n8453), .O(n2936), .CO(n2937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/mVideoTimingGen/add_6/i3  (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .I1(1'b0), .CI(n437), .O(n2938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoTimingGen.v(65)
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i3 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/add_6/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i11  (.I0(\MVideoPostProcess/rVtgRstCnt[10] ), 
            .I1(1'b0), .CI(n2948), .O(n2946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i11 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i10  (.I0(\MVideoPostProcess/rVtgRstCnt[9] ), 
            .I1(1'b0), .CI(n2950), .O(n2947), .CO(n2948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i10 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i9  (.I0(\MVideoPostProcess/rVtgRstCnt[8] ), 
            .I1(1'b0), .CI(n2952), .O(n2949), .CO(n2950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i9 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i8  (.I0(\MVideoPostProcess/rVtgRstCnt[7] ), 
            .I1(1'b0), .CI(n2954), .O(n2951), .CO(n2952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i8 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i7  (.I0(\MVideoPostProcess/rVtgRstCnt[6] ), 
            .I1(1'b0), .CI(n2956), .O(n2953), .CO(n2954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i7 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i6  (.I0(\MVideoPostProcess/rVtgRstCnt[5] ), 
            .I1(1'b0), .CI(n2958), .O(n2955), .CO(n2956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i6 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i5  (.I0(\MVideoPostProcess/rVtgRstCnt[4] ), 
            .I1(1'b0), .CI(n2960), .O(n2957), .CO(n2958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i5 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MVideoPostProcess/add_8/i4  (.I0(\MVideoPostProcess/rVtgRstCnt[3] ), 
            .I1(1'b0), .CI(n332), .O(n2959), .CO(n2960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MVideoPostProcess\MVideoPostProcess.v(175)
    defparam \MVideoPostProcess/add_8/i4 .I0_POLARITY = 1'b1;
    defparam \MVideoPostProcess/add_8/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I1(1'b0), .CI(n2963), .O(n2961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I1(1'b0), .CI(n2965), .O(n2962), .CO(n2963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I1(1'b0), .CI(n2967), .O(n2964), .CO(n2965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I1(1'b0), .CI(n2969), .O(n2966), .CO(n2967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(1'b0), .CI(n2971), .O(n2968), .CO(n2969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4  (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(1'b0), .CI(n211), .O(n2970), .CO(n2971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoController.v(63)
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i10  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I1(1'b0), .CI(n2974), .O(n2972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i9  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(1'b0), .CI(n2976), .O(n2973), .CO(n2974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i8  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(1'b0), .CI(n2978), .O(n2975), .CO(n2976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i7  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(1'b0), .CI(n2980), .O(n2977), .CO(n2978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i6  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I1(1'b0), .CI(n2982), .O(n2979), .CO(n2980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i5  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(1'b0), .CI(n2984), .O(n2981), .CO(n2982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i4  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(1'b0), .CI(n170), .O(n2983), .CO(n2984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i13  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] ), 
            .I1(1'b0), .CI(n2987), .O(n2985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i13 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i12  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .I1(1'b0), .CI(n2989), .O(n2986), .CO(n2987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i12 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i11  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I1(1'b0), .CI(n2991), .O(n2988), .CO(n2989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i11 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i10  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] ), 
            .I1(1'b0), .CI(n2993), .O(n2990), .CO(n2991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i9  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] ), 
            .I1(1'b0), .CI(n2995), .O(n2992), .CO(n2993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i8  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] ), 
            .I1(1'b0), .CI(n2997), .O(n2994), .CO(n2995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i7  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] ), 
            .I1(1'b0), .CI(n2999), .O(n2996), .CO(n2997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i6  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] ), 
            .I1(1'b0), .CI(n3001), .O(n2998), .CO(n2999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i5  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] ), 
            .I1(1'b0), .CI(n3003), .O(n3000), .CO(n3001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i4  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] ), 
            .I1(1'b0), .CI(n3005), .O(n3002), .CO(n3003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/add_49/i3  (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] ), 
            .I1(1'b0), .CI(n125), .O(n3004), .CO(n3005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsi2Decoder.v(270)
    defparam \MCsiRxController/MCsi2Decoder/add_49/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/add_49/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I1(1'b0), .CI(n3008), .O(n3006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(1'b0), .CI(n3010), .O(n3007), .CO(n3008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(1'b0), .CI(n3012), .O(n3009), .CO(n3010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(1'b0), .CI(n3014), .O(n3011), .CO(n3012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I1(1'b0), .CI(n3016), .O(n3013), .CO(n3014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(1'b0), .CI(n3018), .O(n3015), .CO(n3016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(1'b0), .CI(n3020), .O(n3017), .CO(n3018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3  (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(1'b0), .CI(n117), .O(n3019), .CO(n3020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\fifoDualController.v(84)
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/add_15/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i16  (.I0(\la0_probe6[15] ), .I1(1'b0), 
            .CI(n3023), .O(n3021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i16 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i15  (.I0(\la0_probe6[14] ), .I1(1'b0), 
            .CI(n3025), .O(n3022), .CO(n3023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i15 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i14  (.I0(\la0_probe6[13] ), .I1(1'b0), 
            .CI(n3027), .O(n3024), .CO(n3025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i14 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i13  (.I0(\la0_probe6[12] ), .I1(1'b0), 
            .CI(n3029), .O(n3026), .CO(n3027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i13 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i12  (.I0(\la0_probe6[11] ), .I1(1'b0), 
            .CI(n3031), .O(n3028), .CO(n3029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i12 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i11  (.I0(\la0_probe6[10] ), .I1(1'b0), 
            .CI(n3033), .O(n3030), .CO(n3031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i11 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i10  (.I0(\la0_probe6[9] ), .I1(1'b0), 
            .CI(n3035), .O(n3032), .CO(n3033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i10 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i9  (.I0(\la0_probe6[8] ), .I1(1'b0), 
            .CI(n3037), .O(n3034), .CO(n3035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i9 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i8  (.I0(\la0_probe6[7] ), .I1(1'b0), 
            .CI(n3039), .O(n3036), .CO(n3037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i8 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i7  (.I0(\la0_probe6[6] ), .I1(1'b0), 
            .CI(n3041), .O(n3038), .CO(n3039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i7 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i6  (.I0(\la0_probe6[5] ), .I1(1'b0), 
            .CI(n3043), .O(n3040), .CO(n3041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i6 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i5  (.I0(\la0_probe6[4] ), .I1(1'b0), 
            .CI(n3045), .O(n3042), .CO(n3043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i5 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i4  (.I0(\la0_probe6[3] ), .I1(1'b0), 
            .CI(n3047), .O(n3044), .CO(n3045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i4 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i3  (.I0(\la0_probe6[2] ), .I1(1'b0), 
            .CI(n3049), .O(n3046), .CO(n3047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i3 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \MCsiRxController/add_42/i2  (.I0(\la0_probe6[1] ), .I1(\la0_probe6[0] ), 
            .CI(1'b0), .O(n3048), .CO(n3049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\MCsiRxController\MCsiRxController.v(301)
    defparam \MCsiRxController/add_42/i2 .I0_POLARITY = 1'b1;
    defparam \MCsiRxController/add_42/i2 .I1_POLARITY = 1'b1;
    EFX_RAM10 \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo  (.WCLK(oTestPort[17]), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd }), 
            .WDATA({\la0_probe9[1] , \la0_probe9[0] , \la0_probe8[7] , 
            \la0_probe8[6] , \la0_probe8[5] , \la0_probe8[4] , \la0_probe8[3] , 
            \la0_probe8[2] , \la0_probe8[1] , \la0_probe8[0] }), .WADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] }), 
            .RADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] }), 
            .RDATA({\MCsiRxController/MCsi2Decoder/wFtiRd[9] , \MCsiRxController/MCsi2Decoder/wFtiRd[8] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[7] , \MCsiRxController/MCsi2Decoder/wFtiRd[6] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[5] , \MCsiRxController/MCsi2Decoder/wFtiRd[4] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[3] , \MCsiRxController/MCsi2Decoder/wFtiRd[2] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[1] , \MCsiRxController/MCsi2Decoder/wFtiRd[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=10, WRITE_WIDTH=10, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .READ_WIDTH = 10;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 10;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo  (.WCLK(oTestPort[17]), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, \MCsiRxController/MCsi2Decoder/rDphyHsDataLaneVd }), 
            .WDATA({3'b000, \la0_probe3[0] , \la0_probe9[7] , \la0_probe9[6] , 
            \la0_probe9[5] , \la0_probe9[4] , \la0_probe9[3] , \la0_probe9[2] }), 
            .WADDR({\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] }), 
            .RADDR({\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[9] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[8] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[7] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[6] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[5] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[4] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[3] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[2] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[1] , 
            \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rORP[0] }), 
            .RDATA({Open_0, Open_1, Open_2, \MCsiRxController/MCsi2Decoder/wFtiRd[16] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[15] , \MCsiRxController/MCsi2Decoder/wFtiRd[14] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[13] , \MCsiRxController/MCsi2Decoder/wFtiRd[12] , 
            \MCsiRxController/MCsi2Decoder/wFtiRd[11] , \MCsiRxController/MCsi2Decoder/wFtiRd[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=10, WRITE_WIDTH=10, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .READ_WIDTH = 10;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 10;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo  (.WCLK(iSCLK), 
            .RCLK(iSCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({\MCsiRxController/wHsValid , \MCsiRxController/wHsValid }), 
            .WDATA({\MCsiRxController/wHsPixel[15] , \MCsiRxController/wHsPixel[14] , 
            \MCsiRxController/wHsPixel[13] , \MCsiRxController/wHsPixel[12] , 
            \MCsiRxController/wHsPixel[11] , \MCsiRxController/wHsPixel[10] , 
            \MCsiRxController/wHsPixel[9] , \MCsiRxController/wHsPixel[8] , 
            \MCsiRxController/wHsPixel[7] , \MCsiRxController/wHsPixel[6] , 
            \MCsiRxController/wHsPixel[5] , \MCsiRxController/wHsPixel[4] , 
            \MCsiRxController/wHsPixel[3] , \MCsiRxController/wHsPixel[2] , 
            \MCsiRxController/wHsPixel[1] , \MCsiRxController/wHsPixel[0] }), 
            .WADDR({\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] , \MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] }), .RADDR({\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] , 
            \MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] , \MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] }), 
            .RDATA({\wVideoPixel[15] , \wVideoPixel[14] , \wVideoPixel[13] , 
            \wVideoPixel[12] , \wVideoPixel[11] , \wVideoPixel[10] , \wVideoPixel[9] , 
            \wVideoPixel[8] , \wVideoPixel[7] , \wVideoPixel[6] , \wVideoPixel[5] , 
            \wVideoPixel[4] , \wVideoPixel[3] , \wVideoPixel[2] , \wVideoPixel[1] , 
            \wVideoPixel[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=16, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="NONE", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .READ_WIDTH = 16;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WRITE_WIDTH = 16;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WE_POLARITY = 2'b11;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RCLK_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RST_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RESET_RAM = "ASYNC";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RESET_OUTREG = "NONE";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .RE_POLARITY = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .OUTPUT_REG = 1'b1;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .WRITE_MODE = "READ_FIRST";
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MCsiRxController/genblk1[0].mVideoFIFO/USER_FIFO/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram  (.WCLK(1'b0), 
            .RCLK(iBCLK), .WCLKE(1'b0), .RE(1'b1), .RST(1'b0), .WADDREN(1'b0), 
            .RADDREN(1'b1), .WE({2'b00}), .WADDR({10'b0000000000}), .RADDR({\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] , \MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] , 
            \MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] , \MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] , 
            \MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] }), .RDATA({\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] , \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] , 
            \MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=8, WRITE_WIDTH=8, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="NONE", INIT_0=256'h1F24AD230422DC211D201B1F1C1E001D001CAD1B041A3419E71838160115C0D6, INIT_1=256'hC0962856005508481041772F1B2E7C2D082CAD2B042A00290028352701262425, INIT_2=256'h007F00F980FEE0FDE09A01DFD0E0C0D660BA06AFA4A3A4A2619D309CE09A0398, INIT_3=256'h0000000000000000000000000000000000000000000000000000104101E20094, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .READ_WIDTH = 8;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WRITE_WIDTH = 8;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RESET_OUTREG = "NONE";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_0 = 256'h1F24AD230422DC211D201B1F1C1E001D001CAD1B041A3419E71838160115C0D6;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1 = 256'hC0962856005508481041772F1B2E7C2D082CAD2B042A00290028352701262425;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_2 = 256'h007F00F980FEE0FDE09A01DFD0E0C0D660BA06AFA4A3A4A2619D309CE09A0398;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000104101E20094;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .OUTPUT_REG = 1'b1;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/inst_adv7511_config/inst_adv7511_reg/ram .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_SRL8 \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2  (.D(\MVideoPostProcess/mVideoTimingGen/qVrange ), 
            .CLK(iVCLK), .CE(1'b1), .Q(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1 */ ;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .INIT = 8'h0;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_27/i4_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2  (.D(\MVideoPostProcess/mVideoTimingGen/qHrange ), 
            .CLK(iVCLK), .CE(1'b1), .Q(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1 */ ;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .INIT = 8'h0;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .CLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/mVideoTimingGen/dff_11/i4_2 .CE_POLARITY = 1'b1;
    EFX_RAM10 \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[3] , 
            \wVideoPixel[2] , \wVideoPixel[1] , \wVideoPixel[0] }), .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[11:8]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 4;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 4;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[7] , 
            \wVideoPixel[6] , \wVideoPixel[5] , \wVideoPixel[4] }), .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[15:12]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 4;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 4;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[11] , 
            \wVideoPixel[10] , \wVideoPixel[9] , \wVideoPixel[8] }), .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[3:0]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 4;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 4;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo  (.WCLK(iSCLK), 
            .RCLK(iVCLK), .WCLKE(1'b1), .RE(1'b1), .RST(1'b0), .WADDREN(1'b1), 
            .RADDREN(1'b1), .WE({1'b0, wVideoVd}), .WDATA({\wVideoPixel[15] , 
            \wVideoPixel[14] , \wVideoPixel[13] , \wVideoPixel[12] }), 
            .WADDR({\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] , \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] , 
            \MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] }), 
            .RADDR({\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[10] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[9] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[8] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[7] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[6] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[5] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[4] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[3] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[2] , 
            \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[1] , \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rORP[0] }), 
            .RDATA({oAdv7511Data[7:4]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=4, WRITE_WIDTH=4, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .READ_WIDTH = 4;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_WIDTH = 4;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WCLKE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WE_POLARITY = 2'b11;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RCLK_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RST_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RADDREN_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_RAM = "ASYNC";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RESET_OUTREG = "ASYNC";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .RE_POLARITY = 1'b1;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .OUTPUT_REG = 1'b0;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .WRITE_MODE = "READ_UNKNOWN";
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/USER_FIFO_DUAL/fifo .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_LUT4 \edb_top_inst/LUT__3985  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/edb_user_dr[67] ), .I2(\edb_top_inst/la0/crc_data_out[18] ), 
            .I3(\edb_top_inst/edb_user_dr[68] ), .O(\edb_top_inst/n2759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3985 .LUTMASK = 16'h9009;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[2] , \edb_top_inst/la0/la_biu_inst/fifo_dout[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] }), 
            .WADDR({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2  (.D(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_2  (.D(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_2 .CE_POLARITY = 1'b1;
    EFX_SRL8 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2  (.D(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .CLK(oTestPort[17]), .CE(1'b1), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre ), 
            .A({3'b100})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_SRL8, INIT=8'h0, CLK_POLARITY=1'b1, CE_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_SRL8=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .INIT = 8'h0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_2 .CE_POLARITY = 1'b1;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[4] , \edb_top_inst/la0/la_biu_inst/fifo_dout[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[6] , \edb_top_inst/la0/la_biu_inst/fifo_dout[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[8] , \edb_top_inst/la0/la_biu_inst/fifo_dout[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[10] , \edb_top_inst/la0/la_biu_inst/fifo_dout[9] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[12] , \edb_top_inst/la0/la_biu_inst/fifo_dout[11] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[14] , \edb_top_inst/la0/la_biu_inst/fifo_dout[13] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[16] , \edb_top_inst/la0/la_biu_inst/fifo_dout[15] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[18] , \edb_top_inst/la0/la_biu_inst/fifo_dout[17] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[20] , \edb_top_inst/la0/la_biu_inst/fifo_dout[19] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[22] , \edb_top_inst/la0/la_biu_inst/fifo_dout[21] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[24] , \edb_top_inst/la0/la_biu_inst/fifo_dout[23] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[26] , \edb_top_inst/la0/la_biu_inst/fifo_dout[25] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[28] , \edb_top_inst/la0/la_biu_inst/fifo_dout[27] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[30] , \edb_top_inst/la0/la_biu_inst/fifo_dout[29] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$o12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[32] , \edb_top_inst/la0/la_biu_inst/fifo_dout[31] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$p12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[34] , \edb_top_inst/la0/la_biu_inst/fifo_dout[33] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$q12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[36] , \edb_top_inst/la0/la_biu_inst/fifo_dout[35] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$r12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[38] , \edb_top_inst/la0/la_biu_inst/fifo_dout[37] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$s12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[40] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[40] , \edb_top_inst/la0/la_biu_inst/fifo_dout[39] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$t12 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_RAM10 \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1  (.WCLK(oTestPort[17]), 
            .RCLK(oTestPort[17]), .WCLKE(1'b1), .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 ), 
            .RST(1'b0), .WADDREN(1'b1), .RADDREN(1'b1), .WE({1'b0, \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 }), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[42] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[41] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[42] , \edb_top_inst/la0/la_biu_inst/fifo_dout[41] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM10, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=2'b11, WADDREN_POLARITY=1'b1, RADDREN_POLARITY=1'b1, RST_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", RESET_RAM="ASYNC", RESET_OUTREG="ASYNC", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_14=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_15=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_16=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_17=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_18=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_19=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_20=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_21=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_22=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_23=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_24=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_25=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_26=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_27=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM10=TRUE */ ;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WE_POLARITY = 2'b11;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RST_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RADDREN_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RESET_RAM = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RESET_OUTREG = "ASYNC";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .WRITE_MODE = "READ_FIRST";
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$u1 .INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    EFX_LUT4 \edb_top_inst/LUT__3986  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/edb_user_dr[69] ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .I3(\edb_top_inst/edb_user_dr[70] ), .O(\edb_top_inst/n2760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3986 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3987  (.I0(\edb_top_inst/la0/crc_data_out[16] ), 
            .I1(\edb_top_inst/edb_user_dr[66] ), .I2(\edb_top_inst/la0/crc_data_out[23] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n2761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3987 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3988  (.I0(\edb_top_inst/n2758 ), .I1(\edb_top_inst/n2759 ), 
            .I2(\edb_top_inst/n2760 ), .I3(\edb_top_inst/n2761 ), .O(\edb_top_inst/n2762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3988 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3989  (.I0(\edb_top_inst/la0/crc_data_out[24] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .I3(\edb_top_inst/edb_user_dr[81] ), .O(\edb_top_inst/n2763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3989 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3990  (.I0(\edb_top_inst/la0/crc_data_out[25] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/la0/crc_data_out[26] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n2764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3990 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3991  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/edb_user_dr[79] ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n2765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3991 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3992  (.I0(\edb_top_inst/la0/crc_data_out[27] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .I3(\edb_top_inst/edb_user_dr[78] ), .O(\edb_top_inst/n2766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3992 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3993  (.I0(\edb_top_inst/n2763 ), .I1(\edb_top_inst/n2764 ), 
            .I2(\edb_top_inst/n2765 ), .I3(\edb_top_inst/n2766 ), .O(\edb_top_inst/n2767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3993 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3994  (.I0(\edb_top_inst/la0/crc_data_out[0] ), 
            .I1(\edb_top_inst/edb_user_dr[50] ), .I2(\edb_top_inst/la0/crc_data_out[1] ), 
            .I3(\edb_top_inst/edb_user_dr[51] ), .O(\edb_top_inst/n2768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3994 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3995  (.I0(\edb_top_inst/la0/crc_data_out[6] ), 
            .I1(\edb_top_inst/edb_user_dr[56] ), .I2(\edb_top_inst/la0/crc_data_out[15] ), 
            .I3(\edb_top_inst/edb_user_dr[65] ), .O(\edb_top_inst/n2769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3995 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3996  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/edb_user_dr[54] ), .I2(\edb_top_inst/la0/crc_data_out[5] ), 
            .I3(\edb_top_inst/edb_user_dr[55] ), .O(\edb_top_inst/n2770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3996 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3997  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/edb_user_dr[52] ), .I2(\edb_top_inst/la0/crc_data_out[3] ), 
            .I3(\edb_top_inst/edb_user_dr[53] ), .O(\edb_top_inst/n2771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3997 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3998  (.I0(\edb_top_inst/n2768 ), .I1(\edb_top_inst/n2769 ), 
            .I2(\edb_top_inst/n2770 ), .I3(\edb_top_inst/n2771 ), .O(\edb_top_inst/n2772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3998 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3999  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/edb_user_dr[58] ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .I3(\edb_top_inst/edb_user_dr[59] ), .O(\edb_top_inst/n2773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3999 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4000  (.I0(\edb_top_inst/la0/crc_data_out[10] ), 
            .I1(\edb_top_inst/edb_user_dr[60] ), .I2(\edb_top_inst/la0/crc_data_out[11] ), 
            .I3(\edb_top_inst/edb_user_dr[61] ), .O(\edb_top_inst/n2774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4000 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4001  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/edb_user_dr[62] ), .I2(\edb_top_inst/la0/crc_data_out[13] ), 
            .I3(\edb_top_inst/edb_user_dr[63] ), .O(\edb_top_inst/n2775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4001 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4002  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/edb_user_dr[57] ), .I2(\edb_top_inst/la0/crc_data_out[14] ), 
            .I3(\edb_top_inst/edb_user_dr[64] ), .O(\edb_top_inst/n2776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4002 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4003  (.I0(\edb_top_inst/n2773 ), .I1(\edb_top_inst/n2774 ), 
            .I2(\edb_top_inst/n2775 ), .I3(\edb_top_inst/n2776 ), .O(\edb_top_inst/n2777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4003 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4004  (.I0(\edb_top_inst/n2762 ), .I1(\edb_top_inst/n2767 ), 
            .I2(\edb_top_inst/n2772 ), .I3(\edb_top_inst/n2777 ), .O(\edb_top_inst/n2778 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4004 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4005  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(\edb_top_inst/la0/bit_count[3] ), .I2(\edb_top_inst/la0/bit_count[4] ), 
            .I3(\edb_top_inst/la0/bit_count[5] ), .O(\edb_top_inst/n2779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4005 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4006  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/n2779 ), 
            .O(\edb_top_inst/n2780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4006 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4007  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/n2780 ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4007 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4008  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n2782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4008 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4009  (.I0(\edb_top_inst/n2781 ), .I1(\edb_top_inst/n2782 ), 
            .O(\edb_top_inst/n2783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4009 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4010  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/n2778 ), .I2(\edb_top_inst/n2783 ), .O(\edb_top_inst/n2784 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4010 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4011  (.I0(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I1(\edb_top_inst/la0/crc_data_out[0] ), .I2(\edb_top_inst/n2783 ), 
            .O(\edb_top_inst/n2785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4011 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4012  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/n2780 ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n2786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4012 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__4013  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/n2786 ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n2787 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4013 .LUTMASK = 16'h0a0c;
    EFX_LUT4 \edb_top_inst/LUT__4014  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg[1] ), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg[2] ), .I2(\edb_top_inst/debug_hub_inst/module_id_reg[3] ), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg[0] ), .O(\edb_top_inst/n2788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4014 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4015  (.I0(\edb_top_inst/n2785 ), .I1(\edb_top_inst/n2784 ), 
            .I2(\edb_top_inst/n2787 ), .I3(\edb_top_inst/n2788 ), .O(jtag_inst2_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4015 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4016  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[40] ), .O(\edb_top_inst/la0/n1340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4016 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4017  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(jtag_inst2_UPDATE), .I2(\edb_top_inst/n2788 ), .O(\edb_top_inst/n2789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4017 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4018  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n2790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4018 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4019  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .I2(\edb_top_inst/n2790 ), 
            .O(\edb_top_inst/n2791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4019 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4020  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/edb_user_dr[68] ), .I2(\edb_top_inst/edb_user_dr[69] ), 
            .I3(\edb_top_inst/edb_user_dr[79] ), .O(\edb_top_inst/n2792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4020 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4021  (.I0(\edb_top_inst/edb_user_dr[78] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/edb_user_dr[80] ), 
            .O(\edb_top_inst/n2793 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4021 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4022  (.I0(\edb_top_inst/n2789 ), .I1(\edb_top_inst/n2791 ), 
            .I2(\edb_top_inst/n2792 ), .I3(\edb_top_inst/n2793 ), .O(\edb_top_inst/n2794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4022 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4023  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n2794 ), .O(\edb_top_inst/n2795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4023 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4024  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n2795 ), 
            .O(\edb_top_inst/n2796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4024 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4025  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n2797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4025 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4026  (.I0(\edb_top_inst/edb_user_dr[75] ), 
            .I1(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n2798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4026 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4027  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/n2797 ), 
            .I3(\edb_top_inst/n2798 ), .O(\edb_top_inst/n2799 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4027 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4028  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2799 ), 
            .O(\edb_top_inst/la0/n1312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4028 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4029  (.I0(\edb_top_inst/la0/n1312 ), .I1(\edb_top_inst/la0/la_soft_reset_in ), 
            .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4029 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4030  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[41] ), .O(\edb_top_inst/la0/n1341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4030 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4031  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[42] ), .O(\edb_top_inst/la0/n1342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4031 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4032  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n2795 ), 
            .O(\edb_top_inst/n2800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4032 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4033  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2799 ), 
            .O(\edb_top_inst/la0/n1396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4033 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4034  (.I0(\edb_top_inst/n2795 ), .I1(\edb_top_inst/n2799 ), 
            .I2(\edb_top_inst/edb_user_dr[64] ), .I3(\edb_top_inst/edb_user_dr[65] ), 
            .O(\edb_top_inst/la0/n1913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4034 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4035  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/edb_user_dr[63] ), 
            .I3(\edb_top_inst/edb_user_dr[66] ), .O(\edb_top_inst/n2801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4035 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4036  (.I0(\edb_top_inst/n2794 ), .I1(\edb_top_inst/n2799 ), 
            .I2(\edb_top_inst/n2801 ), .O(\edb_top_inst/la0/n1965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4036 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4037  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(\edb_top_inst/la0/address_counter[5] ), .I2(\edb_top_inst/la0/address_counter[6] ), 
            .I3(\edb_top_inst/la0/address_counter[7] ), .O(\edb_top_inst/n2802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4037 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4038  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/address_counter[1] ), .I2(\edb_top_inst/la0/address_counter[2] ), 
            .I3(\edb_top_inst/n2802 ), .O(\edb_top_inst/n2803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4038 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4039  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(\edb_top_inst/la0/address_counter[9] ), .I2(\edb_top_inst/la0/address_counter[10] ), 
            .I3(\edb_top_inst/la0/address_counter[11] ), .O(\edb_top_inst/n2804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4039 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4040  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/la0/address_counter[12] ), .I2(\edb_top_inst/la0/address_counter[13] ), 
            .I3(\edb_top_inst/la0/address_counter[14] ), .O(\edb_top_inst/n2805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4040 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4041  (.I0(\edb_top_inst/n2803 ), .I1(\edb_top_inst/n2804 ), 
            .I2(\edb_top_inst/n2805 ), .O(\edb_top_inst/n2806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4041 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4042  (.I0(\edb_top_inst/n2806 ), .I1(\edb_top_inst/n67 ), 
            .I2(\edb_top_inst/edb_user_dr[45] ), .I3(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4042 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4043  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .I3(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/n2807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4043 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4044  (.I0(\edb_top_inst/n2807 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n2808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4044 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4045  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n2809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4045 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4046  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[6] ), 
            .I3(\edb_top_inst/n2809 ), .O(\edb_top_inst/n2810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4046 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4047  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n2811 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4047 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4048  (.I0(\edb_top_inst/la0/word_count[1] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/la0/word_count[7] ), 
            .I3(\edb_top_inst/la0/word_count[8] ), .O(\edb_top_inst/n2812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4048 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4049  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/n2812 ), .O(\edb_top_inst/n2813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4049 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4050  (.I0(\edb_top_inst/la0/word_count[9] ), 
            .I1(\edb_top_inst/la0/word_count[10] ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .I3(\edb_top_inst/la0/word_count[12] ), .O(\edb_top_inst/n2814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4050 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4051  (.I0(\edb_top_inst/la0/word_count[3] ), 
            .I1(\edb_top_inst/la0/word_count[6] ), .I2(\edb_top_inst/la0/word_count[13] ), 
            .I3(\edb_top_inst/la0/word_count[15] ), .O(\edb_top_inst/n2815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4051 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4052  (.I0(\edb_top_inst/n2813 ), .I1(\edb_top_inst/n2814 ), 
            .I2(\edb_top_inst/n2815 ), .O(\edb_top_inst/n2816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4052 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4053  (.I0(\edb_top_inst/n2810 ), .I1(\edb_top_inst/n2808 ), 
            .I2(\edb_top_inst/n2816 ), .I3(\edb_top_inst/n2811 ), .O(\edb_top_inst/n2817 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5f0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4053 .LUTMASK = 16'h5f0c;
    EFX_LUT4 \edb_top_inst/LUT__4054  (.I0(\edb_top_inst/n2790 ), .I1(\edb_top_inst/n2817 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n2818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4054 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__4055  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n2819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4055 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__4056  (.I0(\edb_top_inst/n2819 ), .I1(\edb_top_inst/la0/bit_count[0] ), 
            .I2(\edb_top_inst/la0/bit_count[1] ), .I3(\edb_top_inst/la0/bit_count[2] ), 
            .O(\edb_top_inst/n2820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbffd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4056 .LUTMASK = 16'hbffd;
    EFX_LUT4 \edb_top_inst/LUT__4057  (.I0(\edb_top_inst/la0/opcode[3] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n2736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4057 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4058  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n2733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4058 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4059  (.I0(\edb_top_inst/n2736 ), .I1(\edb_top_inst/n2733 ), 
            .I2(\edb_top_inst/la0/bit_count[5] ), .I3(\edb_top_inst/la0/bit_count[4] ), 
            .O(\edb_top_inst/n2821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4059 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__4060  (.I0(\edb_top_inst/la0/opcode[1] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n1249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4060 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4061  (.I0(\edb_top_inst/n2819 ), .I1(\edb_top_inst/n1249 ), 
            .O(\edb_top_inst/n2822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4061 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4062  (.I0(\edb_top_inst/n2820 ), .I1(\edb_top_inst/n2821 ), 
            .I2(\edb_top_inst/n2822 ), .I3(\edb_top_inst/la0/bit_count[3] ), 
            .O(\edb_top_inst/n2823 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4062 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__4063  (.I0(\edb_top_inst/n2816 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/n2823 ), 
            .O(\edb_top_inst/n2824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4063 .LUTMASK = 16'hc100;
    EFX_LUT4 \edb_top_inst/LUT__4064  (.I0(\edb_top_inst/n2824 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n2825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4064 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4065  (.I0(\edb_top_inst/edb_user_dr[77] ), 
            .I1(\edb_top_inst/edb_user_dr[78] ), .I2(\edb_top_inst/edb_user_dr[79] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n2826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4065 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__4066  (.I0(\edb_top_inst/n2826 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/n2789 ), .I3(\edb_top_inst/n2790 ), .O(\edb_top_inst/n2827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4066 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4067  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n2827 ), .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4067 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4068  (.I0(\edb_top_inst/n2825 ), .I1(\edb_top_inst/n2818 ), 
            .I2(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4068 .LUTMASK = 16'hf4f4;
    EFX_LUT4 \edb_top_inst/LUT__4069  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n2828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4069 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4070  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/n2823 ), 
            .I3(\edb_top_inst/n2828 ), .O(\edb_top_inst/n2829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4070 .LUTMASK = 16'h9000;
    EFX_LUT4 \edb_top_inst/LUT__4071  (.I0(\edb_top_inst/n2782 ), .I1(\edb_top_inst/n2790 ), 
            .O(\edb_top_inst/n2830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4071 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4072  (.I0(\edb_top_inst/n2829 ), .I1(\edb_top_inst/n2827 ), 
            .I2(\edb_top_inst/n2808 ), .I3(\edb_top_inst/n2830 ), .O(\edb_top_inst/n2831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4072 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4073  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/n2831 ), .O(\edb_top_inst/la0/n2189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4073 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4074  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4074 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4075  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(\edb_top_inst/n2832 ), .I2(\edb_top_inst/n2788 ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4075 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__4076  (.I0(\edb_top_inst/n2833 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/n2828 ), .O(\edb_top_inst/n2834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4076 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__4077  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/n2782 ), .I2(\edb_top_inst/n2834 ), .I3(\edb_top_inst/n2831 ), 
            .O(\edb_top_inst/ceg_net26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4077 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__4078  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/edb_user_dr[29] ), .I2(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_word_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4078 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4079  (.I0(\edb_top_inst/n2816 ), .I1(\edb_top_inst/n2810 ), 
            .O(\edb_top_inst/n2835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4079 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4080  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4080 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4081  (.I0(\edb_top_inst/n2823 ), .I1(\edb_top_inst/n2835 ), 
            .I2(\edb_top_inst/n2836 ), .I3(\edb_top_inst/n2833 ), .O(\edb_top_inst/n2837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4081 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__4082  (.I0(\edb_top_inst/n2816 ), .I1(\edb_top_inst/n2810 ), 
            .I2(\edb_top_inst/n2832 ), .O(\edb_top_inst/n2838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4082 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4083  (.I0(\edb_top_inst/n2788 ), .I1(jtag_inst2_CAPTURE), 
            .O(\edb_top_inst/n2839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4083 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4084  (.I0(\edb_top_inst/n2810 ), .I1(\edb_top_inst/n2816 ), 
            .I2(\edb_top_inst/n2839 ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4084 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__4085  (.I0(\edb_top_inst/n2823 ), .I1(\edb_top_inst/n2838 ), 
            .I2(\edb_top_inst/n2840 ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4085 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4086  (.I0(jtag_inst2_UPDATE), .I1(\edb_top_inst/la0/biu_ready ), 
            .I2(\edb_top_inst/n2839 ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4086 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4087  (.I0(\edb_top_inst/n2842 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/n2827 ), 
            .O(\edb_top_inst/n2843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4087 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4088  (.I0(\edb_top_inst/n2841 ), .I1(\edb_top_inst/n2837 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/n2843 ), 
            .O(\edb_top_inst/n2844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4088 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__4089  (.I0(\edb_top_inst/n2844 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/n2828 ), .I3(\edb_top_inst/n2831 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4089 .LUTMASK = 16'h10ff;
    EFX_LUT4 \edb_top_inst/LUT__4090  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n2845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec07, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4090 .LUTMASK = 16'hec07;
    EFX_LUT4 \edb_top_inst/LUT__4091  (.I0(\edb_top_inst/la0/internal_register_select[10] ), 
            .I1(\edb_top_inst/la0/internal_register_select[11] ), .I2(\edb_top_inst/la0/internal_register_select[12] ), 
            .O(\edb_top_inst/n2846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4091 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4092  (.I0(\edb_top_inst/la0/internal_register_select[1] ), 
            .I1(\edb_top_inst/la0/internal_register_select[2] ), .I2(\edb_top_inst/la0/internal_register_select[4] ), 
            .I3(\edb_top_inst/la0/internal_register_select[5] ), .O(\edb_top_inst/n2847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4092 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4093  (.I0(\edb_top_inst/la0/internal_register_select[6] ), 
            .I1(\edb_top_inst/la0/internal_register_select[7] ), .I2(\edb_top_inst/la0/internal_register_select[8] ), 
            .I3(\edb_top_inst/la0/internal_register_select[9] ), .O(\edb_top_inst/n2848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4093 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4094  (.I0(\edb_top_inst/n2846 ), .I1(\edb_top_inst/n2847 ), 
            .I2(\edb_top_inst/n2848 ), .O(\edb_top_inst/n2849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4094 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4095  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n2849 ), .O(\edb_top_inst/n2850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4095 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4096  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4096 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4097  (.I0(\edb_top_inst/n2849 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n2852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4097 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4098  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n2852 ), .O(\edb_top_inst/n2853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4098 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4099  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I2(\edb_top_inst/n2845 ), .I3(\edb_top_inst/n2851 ), .O(\edb_top_inst/n2854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4099 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__4100  (.I0(\edb_top_inst/n2828 ), .I1(\edb_top_inst/n2823 ), 
            .I2(\edb_top_inst/n2790 ), .I3(\edb_top_inst/n2808 ), .O(\edb_top_inst/n2855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4100 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__4101  (.I0(\edb_top_inst/la0/data_from_biu[0] ), 
            .I1(\edb_top_inst/n2854 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2856 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4101 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4102  (.I0(\edb_top_inst/n2839 ), .I1(\edb_top_inst/n2791 ), 
            .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4102 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__4103  (.I0(\edb_top_inst/la0/data_out_shift_reg[1] ), 
            .I1(\edb_top_inst/n2856 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4103 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4104  (.I0(jtag_inst2_CAPTURE), .I1(jtag_inst2_SHIFT), 
            .I2(\edb_top_inst/n2788 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n2858 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4104 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__4105  (.I0(\edb_top_inst/n2858 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .I2(\edb_top_inst/n2790 ), .I3(\edb_top_inst/n2808 ), .O(\edb_top_inst/ceg_net14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4105 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4106  (.I0(\edb_top_inst/n2780 ), .I1(\edb_top_inst/n2835 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2859 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4106 .LUTMASK = 16'h050c;
    EFX_LUT4 \edb_top_inst/LUT__4107  (.I0(\edb_top_inst/n2859 ), .I1(jtag_inst2_UPDATE), 
            .I2(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n2860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4107 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4108  (.I0(\edb_top_inst/n2860 ), .I1(\edb_top_inst/n2844 ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/la0/module_next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4108 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__4109  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/edb_user_dr[73] ), .I2(\edb_top_inst/n2798 ), 
            .O(\edb_top_inst/n2861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4109 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4110  (.I0(\edb_top_inst/n2861 ), .I1(\edb_top_inst/n2797 ), 
            .O(\edb_top_inst/n2862 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4110 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4111  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2862 ), 
            .O(\edb_top_inst/la0/n5294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4111 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4112  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/n2795 ), .I2(\edb_top_inst/edb_user_dr[65] ), 
            .O(\edb_top_inst/n2863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4112 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4113  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2862 ), 
            .O(\edb_top_inst/la0/n5492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4113 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4114  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2861 ), 
            .O(\edb_top_inst/n2864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4114 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4115  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .O(\edb_top_inst/n2865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4115 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4116  (.I0(\edb_top_inst/n2864 ), .I1(\edb_top_inst/n2865 ), 
            .O(\edb_top_inst/la0/n6947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4116 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4117  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/n2861 ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n2866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4117 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4118  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2866 ), 
            .O(\edb_top_inst/la0/n7907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4118 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4119  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2866 ), 
            .O(\edb_top_inst/la0/n8105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4119 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4120  (.I0(\edb_top_inst/n2798 ), .I1(\edb_top_inst/edb_user_dr[74] ), 
            .O(\edb_top_inst/n2867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4120 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4121  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/n2867 ), .O(\edb_top_inst/n2868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4121 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4122  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2868 ), 
            .O(\edb_top_inst/n2869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4122 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4123  (.I0(\edb_top_inst/n2869 ), .I1(\edb_top_inst/n2797 ), 
            .O(\edb_top_inst/la0/n8741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4123 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4124  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .O(\edb_top_inst/n2870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4124 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4125  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2868 ), 
            .I2(\edb_top_inst/n2870 ), .O(\edb_top_inst/la0/n9645 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4125 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4126  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2868 ), 
            .I2(\edb_top_inst/n2870 ), .O(\edb_top_inst/la0/n9843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4126 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4127  (.I0(\edb_top_inst/n2869 ), .I1(\edb_top_inst/n2865 ), 
            .O(\edb_top_inst/la0/n10527 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4127 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4128  (.I0(\edb_top_inst/n2800 ), .I1(\edb_top_inst/n2868 ), 
            .I2(\edb_top_inst/n2865 ), .O(\edb_top_inst/la0/n10542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4128 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4129  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2868 ), 
            .I2(\edb_top_inst/n2865 ), .O(\edb_top_inst/la0/n10740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4129 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4130  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/n2869 ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/la0/n11368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4130 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4131  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2867 ), 
            .I2(\edb_top_inst/n2797 ), .I3(\edb_top_inst/edb_user_dr[73] ), 
            .O(\edb_top_inst/la0/n12201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4131 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4132  (.I0(\edb_top_inst/n2789 ), .I1(\edb_top_inst/n2791 ), 
            .I2(\edb_top_inst/n2793 ), .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4132 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4133  (.I0(\edb_top_inst/n2806 ), .I1(\edb_top_inst/n1112 ), 
            .I2(\edb_top_inst/edb_user_dr[46] ), .I3(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4133 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4134  (.I0(\edb_top_inst/n2806 ), .I1(\edb_top_inst/n1110 ), 
            .I2(\edb_top_inst/edb_user_dr[47] ), .I3(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4134 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4135  (.I0(\edb_top_inst/n2806 ), .I1(\edb_top_inst/n1108 ), 
            .I2(\edb_top_inst/edb_user_dr[48] ), .I3(\edb_top_inst/n2791 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4135 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4136  (.I0(\edb_top_inst/n1106 ), .I1(\edb_top_inst/edb_user_dr[49] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4136 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4137  (.I0(\edb_top_inst/n1104 ), .I1(\edb_top_inst/edb_user_dr[50] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4137 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4138  (.I0(\edb_top_inst/n1102 ), .I1(\edb_top_inst/edb_user_dr[51] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4138 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4139  (.I0(\edb_top_inst/n1100 ), .I1(\edb_top_inst/edb_user_dr[52] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4139 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4140  (.I0(\edb_top_inst/n1098 ), .I1(\edb_top_inst/edb_user_dr[53] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4140 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4141  (.I0(\edb_top_inst/n1096 ), .I1(\edb_top_inst/edb_user_dr[54] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4141 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4142  (.I0(\edb_top_inst/n1094 ), .I1(\edb_top_inst/edb_user_dr[55] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4142 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4143  (.I0(\edb_top_inst/n1092 ), .I1(\edb_top_inst/edb_user_dr[56] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4143 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4144  (.I0(\edb_top_inst/n1090 ), .I1(\edb_top_inst/edb_user_dr[57] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4144 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4145  (.I0(\edb_top_inst/n1088 ), .I1(\edb_top_inst/edb_user_dr[58] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4145 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4146  (.I0(\edb_top_inst/n1086 ), .I1(\edb_top_inst/edb_user_dr[59] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4146 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4147  (.I0(\edb_top_inst/n1084 ), .I1(\edb_top_inst/la0/address_counter[15] ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2871 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4147 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4148  (.I0(\edb_top_inst/edb_user_dr[60] ), 
            .I1(\edb_top_inst/n2871 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4148 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4149  (.I0(\edb_top_inst/n1082 ), .I1(\edb_top_inst/n1146 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4149 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4150  (.I0(\edb_top_inst/edb_user_dr[61] ), 
            .I1(\edb_top_inst/n2872 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4150 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4151  (.I0(\edb_top_inst/n1080 ), .I1(\edb_top_inst/n1144 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4151 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4152  (.I0(\edb_top_inst/edb_user_dr[62] ), 
            .I1(\edb_top_inst/n2873 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4152 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4153  (.I0(\edb_top_inst/n1078 ), .I1(\edb_top_inst/n1142 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4153 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4154  (.I0(\edb_top_inst/edb_user_dr[63] ), 
            .I1(\edb_top_inst/n2874 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4154 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4155  (.I0(\edb_top_inst/n1076 ), .I1(\edb_top_inst/n1137 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4155 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4156  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/n2875 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4156 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4157  (.I0(\edb_top_inst/n1074 ), .I1(\edb_top_inst/n1135 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4157 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4158  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/n2876 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4158 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4159  (.I0(\edb_top_inst/n1072 ), .I1(\edb_top_inst/n1133 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4159 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4160  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n2877 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4160 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4161  (.I0(\edb_top_inst/n1070 ), .I1(\edb_top_inst/n1131 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4161 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4162  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/n2878 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4162 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4163  (.I0(\edb_top_inst/n1068 ), .I1(\edb_top_inst/n1129 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4163 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4164  (.I0(\edb_top_inst/edb_user_dr[68] ), 
            .I1(\edb_top_inst/n2879 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4164 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4165  (.I0(\edb_top_inst/n1066 ), .I1(\edb_top_inst/n1127 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4165 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4166  (.I0(\edb_top_inst/edb_user_dr[69] ), 
            .I1(\edb_top_inst/n2880 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4166 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4167  (.I0(\edb_top_inst/n1064 ), .I1(\edb_top_inst/n1125 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4167 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4168  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/n2881 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4168 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4169  (.I0(\edb_top_inst/n1062 ), .I1(\edb_top_inst/n1123 ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2882 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4169 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4170  (.I0(\edb_top_inst/edb_user_dr[71] ), 
            .I1(\edb_top_inst/n2882 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_addr_counter[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4170 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4181  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n69 ), 
            .O(\edb_top_inst/la0/n2188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4181 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4182  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n1051 ), 
            .O(\edb_top_inst/la0/n2187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4182 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4183  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n1049 ), 
            .O(\edb_top_inst/la0/n2186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4183 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4184  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n1047 ), 
            .O(\edb_top_inst/la0/n2185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4184 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4185  (.I0(\edb_top_inst/n2831 ), .I1(\edb_top_inst/n1046 ), 
            .O(\edb_top_inst/la0/n2184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4185 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4186  (.I0(\edb_top_inst/edb_user_dr[30] ), 
            .I1(\edb_top_inst/la0/word_count[0] ), .I2(\edb_top_inst/la0/word_count[1] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4186 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__4187  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .O(\edb_top_inst/n2888 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4187 .LUTMASK = 16'he1e1;
    EFX_LUT4 \edb_top_inst/LUT__4188  (.I0(\edb_top_inst/n2888 ), .I1(\edb_top_inst/edb_user_dr[31] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4188 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4189  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n2889 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe01, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4189 .LUTMASK = 16'hfe01;
    EFX_LUT4 \edb_top_inst/LUT__4190  (.I0(\edb_top_inst/n2889 ), .I1(\edb_top_inst/edb_user_dr[32] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4190 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4191  (.I0(\edb_top_inst/edb_user_dr[33] ), 
            .I1(\edb_top_inst/n2809 ), .I2(\edb_top_inst/la0/word_count[4] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4191 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4192  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/n2809 ), .I2(\edb_top_inst/la0/word_count[5] ), 
            .O(\edb_top_inst/n2890 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4192 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4193  (.I0(\edb_top_inst/n2890 ), .I1(\edb_top_inst/edb_user_dr[34] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4193 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4194  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/n2809 ), 
            .I3(\edb_top_inst/la0/word_count[6] ), .O(\edb_top_inst/n2891 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4194 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__4195  (.I0(\edb_top_inst/n2891 ), .I1(\edb_top_inst/edb_user_dr[35] ), 
            .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4195 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4196  (.I0(\edb_top_inst/edb_user_dr[36] ), 
            .I1(\edb_top_inst/n2810 ), .I2(\edb_top_inst/la0/word_count[7] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4196 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4197  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/n2810 ), .I2(\edb_top_inst/la0/word_count[8] ), 
            .O(\edb_top_inst/n2892 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4197 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4198  (.I0(\edb_top_inst/edb_user_dr[37] ), 
            .I1(\edb_top_inst/n2892 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4198 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4199  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/n2810 ), 
            .O(\edb_top_inst/n2893 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4199 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4200  (.I0(\edb_top_inst/edb_user_dr[38] ), 
            .I1(\edb_top_inst/n2893 ), .I2(\edb_top_inst/la0/word_count[9] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4200 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4201  (.I0(\edb_top_inst/la0/word_count[9] ), 
            .I1(\edb_top_inst/n2893 ), .O(\edb_top_inst/n2894 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4201 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4202  (.I0(\edb_top_inst/edb_user_dr[39] ), 
            .I1(\edb_top_inst/n2894 ), .I2(\edb_top_inst/la0/word_count[10] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4202 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4203  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/n2894 ), .O(\edb_top_inst/n2895 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4203 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4204  (.I0(\edb_top_inst/edb_user_dr[40] ), 
            .I1(\edb_top_inst/n2895 ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4204 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4205  (.I0(\edb_top_inst/la0/word_count[11] ), 
            .I1(\edb_top_inst/n2895 ), .O(\edb_top_inst/n2896 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4205 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4206  (.I0(\edb_top_inst/edb_user_dr[41] ), 
            .I1(\edb_top_inst/n2896 ), .I2(\edb_top_inst/la0/word_count[12] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4206 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4207  (.I0(\edb_top_inst/n2893 ), .I1(\edb_top_inst/n2814 ), 
            .O(\edb_top_inst/n2897 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4207 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4208  (.I0(\edb_top_inst/edb_user_dr[42] ), 
            .I1(\edb_top_inst/n2897 ), .I2(\edb_top_inst/la0/word_count[13] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4208 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4209  (.I0(\edb_top_inst/la0/word_count[13] ), 
            .I1(\edb_top_inst/n2897 ), .O(\edb_top_inst/n2898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4209 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4210  (.I0(\edb_top_inst/edb_user_dr[43] ), 
            .I1(\edb_top_inst/n2898 ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4210 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__4211  (.I0(\edb_top_inst/la0/word_count[14] ), 
            .I1(\edb_top_inst/n2898 ), .I2(\edb_top_inst/la0/word_count[15] ), 
            .O(\edb_top_inst/n2899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4211 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__4212  (.I0(\edb_top_inst/edb_user_dr[44] ), 
            .I1(\edb_top_inst/n2899 ), .I2(\edb_top_inst/n2791 ), .O(\edb_top_inst/la0/data_to_word_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4212 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__4213  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2900 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4213 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4214  (.I0(\edb_top_inst/n2851 ), .I1(\edb_top_inst/n2808 ), 
            .I2(\edb_top_inst/n2828 ), .O(\edb_top_inst/n2901 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4214 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4215  (.I0(\edb_top_inst/la0/data_from_biu[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[1] ), .I2(\edb_top_inst/n2900 ), 
            .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4215 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__4216  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4216 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4217  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n2904 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4217 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__4218  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n2903 ), .I2(\edb_top_inst/n2904 ), .O(\edb_top_inst/n2905 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4218 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4219  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n2849 ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .O(\edb_top_inst/n2906 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4219 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4220  (.I0(\edb_top_inst/n2851 ), .I1(\edb_top_inst/n2905 ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4220 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4221  (.I0(\edb_top_inst/n2907 ), .I1(\edb_top_inst/n2902 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[2] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4221 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__4222  (.I0(\edb_top_inst/la0/data_from_biu[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[2] ), .I2(\edb_top_inst/n2900 ), 
            .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4222 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__4223  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n2909 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4223 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4224  (.I0(\edb_top_inst/n2851 ), .I1(\edb_top_inst/n2909 ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2910 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4224 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4225  (.I0(\edb_top_inst/n2910 ), .I1(\edb_top_inst/n2908 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[3] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4225 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__4226  (.I0(\edb_top_inst/la0/data_from_biu[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[3] ), .I2(\edb_top_inst/n2900 ), 
            .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2911 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4226 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4227  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .O(\edb_top_inst/n2912 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d3d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4227 .LUTMASK = 16'h3d3d;
    EFX_LUT4 \edb_top_inst/LUT__4228  (.I0(\edb_top_inst/n2912 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/n2900 ), .O(\edb_top_inst/n2913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4228 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4229  (.I0(\edb_top_inst/n2913 ), .I1(\edb_top_inst/n2911 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[4] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf011, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4229 .LUTMASK = 16'hf011;
    EFX_LUT4 \edb_top_inst/LUT__4230  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[4] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4230 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4231  (.I0(\edb_top_inst/la0/data_from_biu[4] ), 
            .I1(\edb_top_inst/n2914 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2915 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4231 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4232  (.I0(\edb_top_inst/n2915 ), .I1(\edb_top_inst/la0/data_out_shift_reg[5] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4232 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4233  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[5] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2916 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4233 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4234  (.I0(\edb_top_inst/la0/data_from_biu[5] ), 
            .I1(\edb_top_inst/n2916 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2917 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4234 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4235  (.I0(\edb_top_inst/n2917 ), .I1(\edb_top_inst/la0/data_out_shift_reg[6] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4235 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4236  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[6] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2918 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4236 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4237  (.I0(\edb_top_inst/n2918 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[6] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2919 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4237 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4238  (.I0(\edb_top_inst/n2919 ), .I1(\edb_top_inst/la0/data_out_shift_reg[7] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4238 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4239  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[7] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2920 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4239 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4240  (.I0(\edb_top_inst/n2920 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[7] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2921 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4240 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4241  (.I0(\edb_top_inst/n2921 ), .I1(\edb_top_inst/la0/data_out_shift_reg[8] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4241 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4242  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2922 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4242 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4243  (.I0(\edb_top_inst/n2922 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[8] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2923 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4243 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4244  (.I0(\edb_top_inst/n2923 ), .I1(\edb_top_inst/la0/data_out_shift_reg[9] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4244 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4245  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2924 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4245 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4246  (.I0(\edb_top_inst/la0/la_trig_mask[9] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[9] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2925 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4246 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4247  (.I0(\edb_top_inst/n2924 ), .I1(\edb_top_inst/n2925 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[10] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4247 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4248  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[10] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2926 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4248 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4249  (.I0(\edb_top_inst/la0/data_from_biu[10] ), 
            .I1(\edb_top_inst/n2926 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2927 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4249 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4250  (.I0(\edb_top_inst/n2927 ), .I1(\edb_top_inst/la0/data_out_shift_reg[11] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4250 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4251  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[11] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2928 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4251 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4252  (.I0(\edb_top_inst/n2928 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[11] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2929 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4252 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4253  (.I0(\edb_top_inst/n2929 ), .I1(\edb_top_inst/la0/data_out_shift_reg[12] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4253 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4254  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[12] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2930 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4254 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4255  (.I0(\edb_top_inst/n2930 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[12] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2931 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4255 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4256  (.I0(\edb_top_inst/n2931 ), .I1(\edb_top_inst/la0/data_out_shift_reg[13] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4256 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4257  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[13] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2932 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4257 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4258  (.I0(\edb_top_inst/la0/data_from_biu[13] ), 
            .I1(\edb_top_inst/n2932 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2933 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4258 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4259  (.I0(\edb_top_inst/n2933 ), .I1(\edb_top_inst/la0/data_out_shift_reg[14] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4259 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4260  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[14] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2934 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4260 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4261  (.I0(\edb_top_inst/n2934 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[14] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2935 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4261 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4262  (.I0(\edb_top_inst/n2935 ), .I1(\edb_top_inst/la0/data_out_shift_reg[15] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4262 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4263  (.I0(\edb_top_inst/la0/la_sample_cnt[12] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[15] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2936 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4263 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4264  (.I0(\edb_top_inst/n2936 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[15] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2937 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4264 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4265  (.I0(\edb_top_inst/n2937 ), .I1(\edb_top_inst/la0/data_out_shift_reg[16] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4265 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4266  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[16] ), .I2(\edb_top_inst/n2852 ), 
            .O(\edb_top_inst/n2938 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4266 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4267  (.I0(\edb_top_inst/la0/data_from_biu[16] ), 
            .I1(\edb_top_inst/n2938 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2939 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4267 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4268  (.I0(\edb_top_inst/n2939 ), .I1(\edb_top_inst/la0/data_out_shift_reg[17] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4268 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4269  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[17] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/n2849 ), .O(\edb_top_inst/n2940 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4269 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4270  (.I0(\edb_top_inst/la0/data_from_biu[17] ), 
            .I1(\edb_top_inst/n2940 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2941 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4270 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4271  (.I0(\edb_top_inst/n2941 ), .I1(\edb_top_inst/la0/data_out_shift_reg[18] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4271 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4272  (.I0(\edb_top_inst/n2850 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[18] ), .O(\edb_top_inst/n2942 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4272 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4273  (.I0(\edb_top_inst/la0/data_from_biu[18] ), 
            .I1(\edb_top_inst/n2942 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2943 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4273 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4274  (.I0(\edb_top_inst/n2943 ), .I1(\edb_top_inst/la0/data_out_shift_reg[19] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4274 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4275  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[19] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/n2849 ), .O(\edb_top_inst/n2944 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4275 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4276  (.I0(\edb_top_inst/la0/data_from_biu[19] ), 
            .I1(\edb_top_inst/n2944 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2945 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4276 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4277  (.I0(\edb_top_inst/n2945 ), .I1(\edb_top_inst/la0/data_out_shift_reg[20] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4277 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4278  (.I0(\edb_top_inst/la0/la_trig_mask[20] ), 
            .I1(\edb_top_inst/la0/la_run_trig ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2946 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4278 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4279  (.I0(\edb_top_inst/n2946 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[20] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4279 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4280  (.I0(\edb_top_inst/n2947 ), .I1(\edb_top_inst/la0/data_out_shift_reg[21] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4280 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4281  (.I0(\edb_top_inst/la0/la_trig_mask[21] ), 
            .I1(\edb_top_inst/la0/la_run_trig_imdt ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2948 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4281 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4282  (.I0(\edb_top_inst/la0/data_from_biu[21] ), 
            .I1(\edb_top_inst/n2948 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2949 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4282 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4283  (.I0(\edb_top_inst/n2949 ), .I1(\edb_top_inst/la0/data_out_shift_reg[22] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4283 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4284  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2950 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4284 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4285  (.I0(\edb_top_inst/la0/la_trig_mask[22] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[22] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2951 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4285 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4286  (.I0(\edb_top_inst/n2950 ), .I1(\edb_top_inst/n2951 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[23] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4286 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4287  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[23] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2952 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4287 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4288  (.I0(\edb_top_inst/la0/data_from_biu[23] ), 
            .I1(\edb_top_inst/n2952 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2953 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4288 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4289  (.I0(\edb_top_inst/n2953 ), .I1(\edb_top_inst/la0/data_out_shift_reg[24] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4289 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4290  (.I0(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[24] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2954 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4290 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4291  (.I0(\edb_top_inst/n2954 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[24] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2955 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4291 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4292  (.I0(\edb_top_inst/n2955 ), .I1(\edb_top_inst/la0/data_out_shift_reg[25] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4292 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4293  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[25] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2956 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4293 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4294  (.I0(\edb_top_inst/n2956 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[25] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2957 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4294 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4295  (.I0(\edb_top_inst/n2957 ), .I1(\edb_top_inst/la0/data_out_shift_reg[26] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4295 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4296  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[26] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2958 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4296 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4297  (.I0(\edb_top_inst/n2958 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[26] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4297 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4298  (.I0(\edb_top_inst/n2959 ), .I1(\edb_top_inst/la0/data_out_shift_reg[27] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4298 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4299  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[27] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4299 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4300  (.I0(\edb_top_inst/la0/data_from_biu[27] ), 
            .I1(\edb_top_inst/n2960 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2961 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4300 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4301  (.I0(\edb_top_inst/n2961 ), .I1(\edb_top_inst/la0/data_out_shift_reg[28] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4301 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4302  (.I0(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[28] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2962 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4302 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4303  (.I0(\edb_top_inst/la0/data_from_biu[28] ), 
            .I1(\edb_top_inst/n2962 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2963 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4303 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4304  (.I0(\edb_top_inst/n2963 ), .I1(\edb_top_inst/la0/data_out_shift_reg[29] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4304 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4305  (.I0(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[29] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2964 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4305 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4306  (.I0(\edb_top_inst/la0/data_from_biu[29] ), 
            .I1(\edb_top_inst/n2964 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4306 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4307  (.I0(\edb_top_inst/n2965 ), .I1(\edb_top_inst/la0/data_out_shift_reg[30] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4307 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4308  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[30] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4308 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4309  (.I0(\edb_top_inst/n2966 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[30] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2967 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4309 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4310  (.I0(\edb_top_inst/n2967 ), .I1(\edb_top_inst/la0/data_out_shift_reg[31] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4310 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4311  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[31] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2968 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4311 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4312  (.I0(\edb_top_inst/la0/data_from_biu[31] ), 
            .I1(\edb_top_inst/n2968 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2969 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4312 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4313  (.I0(\edb_top_inst/n2969 ), .I1(\edb_top_inst/la0/data_out_shift_reg[32] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4313 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4314  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4314 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4315  (.I0(\edb_top_inst/la0/la_trig_mask[32] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[32] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2971 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4315 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4316  (.I0(\edb_top_inst/n2970 ), .I1(\edb_top_inst/n2971 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[33] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4316 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4317  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4317 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4318  (.I0(\edb_top_inst/la0/la_trig_mask[33] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[33] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2973 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4318 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4319  (.I0(\edb_top_inst/n2972 ), .I1(\edb_top_inst/n2973 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[34] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4319 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4320  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[34] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4320 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4321  (.I0(\edb_top_inst/la0/data_from_biu[34] ), 
            .I1(\edb_top_inst/n2974 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2975 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4321 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4322  (.I0(\edb_top_inst/n2975 ), .I1(\edb_top_inst/la0/data_out_shift_reg[35] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4322 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4323  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2976 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4323 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4324  (.I0(\edb_top_inst/la0/la_trig_mask[35] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[35] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2977 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4324 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4325  (.I0(\edb_top_inst/n2976 ), .I1(\edb_top_inst/n2977 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[36] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4325 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4326  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[36] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2978 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4326 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4327  (.I0(\edb_top_inst/la0/data_from_biu[36] ), 
            .I1(\edb_top_inst/n2978 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2979 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4327 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4328  (.I0(\edb_top_inst/n2979 ), .I1(\edb_top_inst/la0/data_out_shift_reg[37] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4328 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4329  (.I0(\edb_top_inst/la0/la_trig_pos[14] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[37] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2980 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4329 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4330  (.I0(\edb_top_inst/n2980 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[37] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2981 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4330 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4331  (.I0(\edb_top_inst/n2981 ), .I1(\edb_top_inst/la0/data_out_shift_reg[38] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4331 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4332  (.I0(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[38] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2982 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4332 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4333  (.I0(\edb_top_inst/n2982 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[38] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2983 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4333 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4334  (.I0(\edb_top_inst/n2983 ), .I1(\edb_top_inst/la0/data_out_shift_reg[39] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4334 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4335  (.I0(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[39] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2984 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4335 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4336  (.I0(\edb_top_inst/n2984 ), .I1(\edb_top_inst/n2849 ), 
            .I2(\edb_top_inst/la0/data_from_biu[39] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2985 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4336 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4337  (.I0(\edb_top_inst/n2985 ), .I1(\edb_top_inst/la0/data_out_shift_reg[40] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4337 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4338  (.I0(\edb_top_inst/la0/la_trig_mask[40] ), 
            .I1(\edb_top_inst/la0/la_trig_pattern[0] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2986 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4338 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__4339  (.I0(\edb_top_inst/la0/data_from_biu[40] ), 
            .I1(\edb_top_inst/n2986 ), .I2(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4339 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4340  (.I0(\edb_top_inst/n2987 ), .I1(\edb_top_inst/la0/data_out_shift_reg[41] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4340 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__4341  (.I0(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[41] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2988 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4341 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4342  (.I0(\edb_top_inst/n2988 ), .I1(\edb_top_inst/n2906 ), 
            .I2(\edb_top_inst/la0/data_from_biu[41] ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2989 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4342 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__4343  (.I0(\edb_top_inst/n2989 ), .I1(\edb_top_inst/la0/data_out_shift_reg[42] ), 
            .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4343 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4344  (.I0(\edb_top_inst/la0/la_capture_pattern[0] ), 
            .I1(\edb_top_inst/n2901 ), .I2(\edb_top_inst/n2852 ), .I3(\edb_top_inst/n2855 ), 
            .O(\edb_top_inst/n2990 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4344 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4345  (.I0(\edb_top_inst/la0/la_trig_mask[42] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/la0/data_from_biu[42] ), 
            .I3(\edb_top_inst/n2855 ), .O(\edb_top_inst/n2991 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4345 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__4346  (.I0(\edb_top_inst/n2990 ), .I1(\edb_top_inst/n2991 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[43] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4346 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__4347  (.I0(\edb_top_inst/la0/la_capture_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[43] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2850 ), .O(\edb_top_inst/n2992 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4347 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4348  (.I0(\edb_top_inst/n2855 ), .I1(\edb_top_inst/n2992 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[44] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4348 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4349  (.I0(\edb_top_inst/n2855 ), .I1(\edb_top_inst/n2853 ), 
            .O(\edb_top_inst/n2993 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4349 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4350  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[44] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[45] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4350 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4351  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[45] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2994 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4351 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4352  (.I0(\edb_top_inst/la0/data_out_shift_reg[46] ), 
            .I1(\edb_top_inst/n2994 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4352 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4353  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[46] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2995 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4353 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4354  (.I0(\edb_top_inst/la0/data_out_shift_reg[47] ), 
            .I1(\edb_top_inst/n2995 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4354 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4355  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[47] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n2996 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4355 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4356  (.I0(\edb_top_inst/la0/data_out_shift_reg[48] ), 
            .I1(\edb_top_inst/n2996 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4356 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4357  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[48] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[49] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4357 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4358  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[49] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2997 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4358 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4359  (.I0(\edb_top_inst/la0/data_out_shift_reg[50] ), 
            .I1(\edb_top_inst/n2997 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4359 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4360  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[50] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[51] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4360 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4361  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[51] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2998 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4361 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4362  (.I0(\edb_top_inst/la0/data_out_shift_reg[52] ), 
            .I1(\edb_top_inst/n2998 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4362 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4363  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[52] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[53] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4363 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4364  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[53] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n2999 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4364 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4365  (.I0(\edb_top_inst/la0/data_out_shift_reg[54] ), 
            .I1(\edb_top_inst/n2999 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4365 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4366  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[54] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n3000 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4366 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4367  (.I0(\edb_top_inst/la0/data_out_shift_reg[55] ), 
            .I1(\edb_top_inst/n3000 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4367 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4368  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[55] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2849 ), .O(\edb_top_inst/n3001 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4368 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4369  (.I0(\edb_top_inst/la0/data_out_shift_reg[56] ), 
            .I1(\edb_top_inst/n3001 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4369 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4370  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[56] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n3002 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4370 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4371  (.I0(\edb_top_inst/la0/data_out_shift_reg[57] ), 
            .I1(\edb_top_inst/n3002 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4371 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4372  (.I0(\edb_top_inst/n2993 ), .I1(\edb_top_inst/la0/la_trig_mask[57] ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[58] ), .I3(\edb_top_inst/n2857 ), 
            .O(\edb_top_inst/la0/n2409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf088, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4372 .LUTMASK = 16'hf088;
    EFX_LUT4 \edb_top_inst/LUT__4373  (.I0(\edb_top_inst/n2853 ), .I1(\edb_top_inst/la0/la_trig_mask[58] ), 
            .I2(\edb_top_inst/n2906 ), .I3(\edb_top_inst/n2901 ), .O(\edb_top_inst/n3003 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4373 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4374  (.I0(\edb_top_inst/la0/data_out_shift_reg[59] ), 
            .I1(\edb_top_inst/n3003 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4374 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4375  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[59] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2849 ), .O(\edb_top_inst/n3004 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4375 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4376  (.I0(\edb_top_inst/la0/data_out_shift_reg[60] ), 
            .I1(\edb_top_inst/n3004 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4376 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4377  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[60] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n3005 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4377 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4378  (.I0(\edb_top_inst/la0/data_out_shift_reg[61] ), 
            .I1(\edb_top_inst/n3005 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4378 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4379  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[61] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n3006 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4379 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4380  (.I0(\edb_top_inst/la0/data_out_shift_reg[62] ), 
            .I1(\edb_top_inst/n3006 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4380 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4381  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[62] ), .I2(\edb_top_inst/n2901 ), 
            .I3(\edb_top_inst/n2852 ), .O(\edb_top_inst/n3007 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4381 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4382  (.I0(\edb_top_inst/la0/data_out_shift_reg[63] ), 
            .I1(\edb_top_inst/n3007 ), .I2(\edb_top_inst/n2857 ), .O(\edb_top_inst/la0/n2404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4382 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__4383  (.I0(\edb_top_inst/la0/la_trig_mask[63] ), 
            .I1(\edb_top_inst/n2853 ), .I2(\edb_top_inst/n2906 ), .O(\edb_top_inst/n3008 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4383 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4384  (.I0(\edb_top_inst/n2857 ), .I1(\edb_top_inst/n3008 ), 
            .I2(\edb_top_inst/n2901 ), .O(\edb_top_inst/la0/n2403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4384 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4385  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/biu_ready ), .I2(jtag_inst2_UPDATE), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n3009 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f57, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4385 .LUTMASK = 16'h0f57;
    EFX_LUT4 \edb_top_inst/LUT__4386  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n2839 ), .I2(\edb_top_inst/n2835 ), .I3(\edb_top_inst/n2811 ), 
            .O(\edb_top_inst/n3010 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4386 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4387  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/n3009 ), .I2(\edb_top_inst/n3010 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n3011 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4387 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__4388  (.I0(\edb_top_inst/n2811 ), .I1(jtag_inst2_UPDATE), 
            .I2(\edb_top_inst/n2782 ), .I3(\edb_top_inst/n3011 ), .O(\edb_top_inst/la0/module_next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4388 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__4389  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/n2823 ), 
            .I3(\edb_top_inst/n2828 ), .O(\edb_top_inst/n3012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4389 .LUTMASK = 16'hb200;
    EFX_LUT4 \edb_top_inst/LUT__4390  (.I0(\edb_top_inst/n2830 ), .I1(\edb_top_inst/n3012 ), 
            .I2(\edb_top_inst/n2828 ), .I3(\edb_top_inst/n2835 ), .O(\edb_top_inst/n3013 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h30fa, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4390 .LUTMASK = 16'h30fa;
    EFX_LUT4 \edb_top_inst/LUT__4391  (.I0(\edb_top_inst/n2808 ), .I1(\edb_top_inst/n3013 ), 
            .I2(\edb_top_inst/n2811 ), .I3(jtag_inst2_UPDATE), .O(\edb_top_inst/la0/module_next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4391 .LUTMASK = 16'he0ee;
    EFX_LUT4 \edb_top_inst/LUT__4392  (.I0(\edb_top_inst/n2790 ), .I1(\edb_top_inst/n2835 ), 
            .I2(\edb_top_inst/n2782 ), .O(\edb_top_inst/n3014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4392 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4393  (.I0(\edb_top_inst/n2835 ), .I1(\edb_top_inst/n2829 ), 
            .I2(\edb_top_inst/n3014 ), .I3(jtag_inst2_UPDATE), .O(\edb_top_inst/la0/module_next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4393 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__4394  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[1] ), .O(\edb_top_inst/la0/axi_crc_i/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4394 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4395  (.I0(\edb_top_inst/n2811 ), .I1(\edb_top_inst/n2782 ), 
            .I2(\edb_top_inst/la0/op_reg_en ), .I3(\edb_top_inst/n2834 ), 
            .O(\edb_top_inst/ceg_net221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4395 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4396  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[2] ), .O(\edb_top_inst/la0/axi_crc_i/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4396 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4397  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[3] ), .O(\edb_top_inst/la0/axi_crc_i/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4397 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4398  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[4] ), .O(\edb_top_inst/la0/axi_crc_i/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4398 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4399  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[5] ), .O(\edb_top_inst/la0/axi_crc_i/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4399 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4400  (.I0(jtag_inst2_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/crc_data_out[0] ), 
            .O(\edb_top_inst/n3015 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4400 .LUTMASK = 16'hac53;
    EFX_LUT4 \edb_top_inst/LUT__4401  (.I0(\edb_top_inst/n3015 ), .I1(\edb_top_inst/n2834 ), 
            .O(\edb_top_inst/n3016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4401 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4402  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[6] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4402 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4403  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[7] ), .O(\edb_top_inst/la0/axi_crc_i/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4403 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4404  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[8] ), .O(\edb_top_inst/la0/axi_crc_i/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4404 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4405  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4405 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4406  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[10] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4406 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4407  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[11] ), .O(\edb_top_inst/la0/axi_crc_i/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4407 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4408  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[12] ), .O(\edb_top_inst/la0/axi_crc_i/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4408 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4409  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[13] ), .O(\edb_top_inst/la0/axi_crc_i/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4409 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4410  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[14] ), .O(\edb_top_inst/la0/axi_crc_i/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4410 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4411  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[15] ), .O(\edb_top_inst/la0/axi_crc_i/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4411 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4412  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[16] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4412 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4413  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[17] ), .O(\edb_top_inst/la0/axi_crc_i/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4413 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4414  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[18] ), .O(\edb_top_inst/la0/axi_crc_i/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4414 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4415  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[19] ), .O(\edb_top_inst/la0/axi_crc_i/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4415 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4416  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4416 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4417  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[21] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4417 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4418  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4418 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4419  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[23] ), .O(\edb_top_inst/la0/axi_crc_i/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4419 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4420  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[24] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4420 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4421  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[25] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4421 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4422  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[26] ), .O(\edb_top_inst/la0/axi_crc_i/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4422 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4423  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[27] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4423 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4424  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4424 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4425  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[29] ), .O(\edb_top_inst/la0/axi_crc_i/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4425 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4426  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4426 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4427  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .O(\edb_top_inst/la0/axi_crc_i/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbebe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4427 .LUTMASK = 16'hbebe;
    EFX_LUT4 \edb_top_inst/LUT__4428  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n3016 ), .O(\edb_top_inst/la0/axi_crc_i/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4428 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4429  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/n2796 ), 
            .I3(\edb_top_inst/n2798 ), .O(\edb_top_inst/n3017 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4429 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4430  (.I0(\edb_top_inst/n3017 ), .I1(\edb_top_inst/n2870 ), 
            .O(\edb_top_inst/la0/n2766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4430 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4431  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4431 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4432  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4432 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4433  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4433 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4434  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4434 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4435  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4435 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4436  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3019 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4436 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4437  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4437 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4438  (.I0(\edb_top_inst/n3019 ), .I1(\edb_top_inst/n3018 ), 
            .I2(\edb_top_inst/n3020 ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4438 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4439  (.I0(\edb_top_inst/n3017 ), .I1(\edb_top_inst/n2865 ), 
            .O(\edb_top_inst/la0/n3599 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4439 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4440  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4440 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4441  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4441 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4442  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4442 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4443  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4443 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4444  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3021 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4444 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4445  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4445 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4446  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3023 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4446 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4447  (.I0(\edb_top_inst/n3022 ), .I1(\edb_top_inst/n3021 ), 
            .I2(\edb_top_inst/n3023 ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4447 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4448  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/n3017 ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/la0/n4432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4448 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4449  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4449 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4450  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4450 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4451  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4451 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4452  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4452 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4453  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3024 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4453 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4454  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3025 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4454 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4455  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3026 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4455 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4456  (.I0(\edb_top_inst/n3025 ), .I1(\edb_top_inst/n3024 ), 
            .I2(\edb_top_inst/n3026 ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4456 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4457  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2862 ), 
            .O(\edb_top_inst/la0/n5279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4457 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4458  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4458 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4459  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4459 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4460  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b22, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4460 .LUTMASK = 16'h2b22;
    EFX_LUT4 \edb_top_inst/LUT__4461  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ff6, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4461 .LUTMASK = 16'h6ff6;
    EFX_LUT4 \edb_top_inst/LUT__4462  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4462 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4463  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n3027 ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3028 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4463 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4464  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3029 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4464 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4465  (.I0(\edb_top_inst/n3027 ), .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n3029 ), .O(\edb_top_inst/n3030 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4c70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4465 .LUTMASK = 16'h4c70;
    EFX_LUT4 \edb_top_inst/LUT__4466  (.I0(\edb_top_inst/n3030 ), .I1(\edb_top_inst/n3028 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4466 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4467  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4467 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4468  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4468 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4469  (.I0(\edb_top_inst/n2864 ), .I1(\edb_top_inst/n2870 ), 
            .O(\edb_top_inst/la0/n6114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4469 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4470  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4470 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4471  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4471 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4472  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4472 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4473  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4473 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4474  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3031 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4474 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4475  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3032 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4475 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4476  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4476 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4477  (.I0(\edb_top_inst/n3032 ), .I1(\edb_top_inst/n3031 ), 
            .I2(\edb_top_inst/n3033 ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4477 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4478  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4478 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4479  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4479 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4480  (.I0(\edb_top_inst/la0/GEN_PROBE[5].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4480 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4481  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4481 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4482  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3034 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4482 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4483  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3035 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4483 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4484  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3036 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4484 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4485  (.I0(\edb_top_inst/n3035 ), .I1(\edb_top_inst/n3034 ), 
            .I2(\edb_top_inst/n3036 ), .I3(\edb_top_inst/la0/GEN_PROBE[5].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4485 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4486  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/n2866 ), 
            .O(\edb_top_inst/la0/n7892 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4486 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4487  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4487 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4488  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4488 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4489  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n3037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4489 .LUTMASK = 16'h8eaf;
    EFX_LUT4 \edb_top_inst/LUT__4490  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), .O(\edb_top_inst/n3038 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4490 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4491  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3039 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4491 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4492  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), .O(\edb_top_inst/n3040 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4492 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4493  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), .O(\edb_top_inst/n3041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4493 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4494  (.I0(\edb_top_inst/n3039 ), .I1(\edb_top_inst/n3038 ), 
            .I2(\edb_top_inst/n3040 ), .I3(\edb_top_inst/n3041 ), .O(\edb_top_inst/n3042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4494 .LUTMASK = 16'hd000;
    EFX_LUT4 \edb_top_inst/LUT__4495  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4495 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4496  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n3044 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4496 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4497  (.I0(\edb_top_inst/n3043 ), .I1(\edb_top_inst/n3040 ), 
            .I2(\edb_top_inst/n3044 ), .O(\edb_top_inst/n3045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4497 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4498  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), .O(\edb_top_inst/n3046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4498 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4499  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3047 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4499 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4500  (.I0(\edb_top_inst/n3042 ), .I1(\edb_top_inst/n3045 ), 
            .I2(\edb_top_inst/n3046 ), .I3(\edb_top_inst/n3047 ), .O(\edb_top_inst/n3048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4500 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__4501  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), .O(\edb_top_inst/n3049 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4501 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4502  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/n3050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4502 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4503  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n3051 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4503 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4504  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), .I2(\edb_top_inst/n3050 ), 
            .I3(\edb_top_inst/n3051 ), .O(\edb_top_inst/n3052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4504 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__4505  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), .O(\edb_top_inst/n3053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4505 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4506  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n3054 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4506 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4507  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), .I2(\edb_top_inst/n3054 ), 
            .O(\edb_top_inst/n3055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4507 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4508  (.I0(\edb_top_inst/n3053 ), .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/n3055 ), .O(\edb_top_inst/n3056 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4508 .LUTMASK = 16'hb200;
    EFX_LUT4 \edb_top_inst/LUT__4509  (.I0(\edb_top_inst/n3048 ), .I1(\edb_top_inst/n3049 ), 
            .I2(\edb_top_inst/n3052 ), .I3(\edb_top_inst/n3056 ), .O(\edb_top_inst/n3057 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4509 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__4510  (.I0(\edb_top_inst/n3037 ), .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), .I3(\edb_top_inst/n3057 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4510 .LUTMASK = 16'h00b2;
    EFX_LUT4 \edb_top_inst/LUT__4511  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), .O(\edb_top_inst/n3058 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4511 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4512  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[0] ), .I2(\edb_top_inst/n3052 ), 
            .I3(\edb_top_inst/n3058 ), .O(\edb_top_inst/n3059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4512 .LUTMASK = 16'hd000;
    EFX_LUT4 \edb_top_inst/LUT__4513  (.I0(\edb_top_inst/n3038 ), .I1(\edb_top_inst/n3039 ), 
            .I2(\edb_top_inst/n3043 ), .I3(\edb_top_inst/n3044 ), .O(\edb_top_inst/n3060 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4513 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4514  (.I0(\edb_top_inst/n3049 ), .I1(\edb_top_inst/n3047 ), 
            .I2(\edb_top_inst/n3046 ), .I3(\edb_top_inst/n3053 ), .O(\edb_top_inst/n3061 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4514 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4515  (.I0(\edb_top_inst/n3055 ), .I1(\edb_top_inst/n3060 ), 
            .I2(\edb_top_inst/n3061 ), .O(\edb_top_inst/n3062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4515 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4516  (.I0(\edb_top_inst/n3059 ), .I1(\edb_top_inst/n3062 ), 
            .I2(\edb_top_inst/n3040 ), .I3(\edb_top_inst/n3041 ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/equal_9/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4516 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4517  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .O(\edb_top_inst/n3063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4517 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4518  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n3064 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4518 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4519  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n3065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4519 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4520  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .O(\edb_top_inst/n3066 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4520 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4521  (.I0(\edb_top_inst/n3063 ), .I1(\edb_top_inst/n3064 ), 
            .I2(\edb_top_inst/n3065 ), .I3(\edb_top_inst/n3066 ), .O(\edb_top_inst/n3067 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4521 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4522  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .O(\edb_top_inst/n3068 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4522 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4523  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .O(\edb_top_inst/n3069 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4523 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4524  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .O(\edb_top_inst/n3070 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4524 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4525  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n3071 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4525 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4526  (.I0(\edb_top_inst/n3068 ), .I1(\edb_top_inst/n3069 ), 
            .I2(\edb_top_inst/n3070 ), .I3(\edb_top_inst/n3071 ), .O(\edb_top_inst/n3072 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4526 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4527  (.I0(\edb_top_inst/n3067 ), .I1(\edb_top_inst/n3072 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/n3073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4527 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__4528  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .I3(\edb_top_inst/n3073 ), .O(\edb_top_inst/n3074 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc513, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4528 .LUTMASK = 16'hc513;
    EFX_LUT4 \edb_top_inst/LUT__4529  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3075 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4529 .LUTMASK = 16'hccca;
    EFX_LUT4 \edb_top_inst/LUT__4530  (.I0(\edb_top_inst/n3075 ), .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/n3074 ), .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4530 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4531  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4531 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4532  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4532 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4533  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4533 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4534  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4534 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4535  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4535 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4536  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4536 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4537  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4537 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4538  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4538 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4539  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4539 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4540  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4540 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4541  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4541 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4542  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4542 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4543  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4543 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4544  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4544 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4545  (.I0(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4545 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4546  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4546 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4547  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4547 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4548  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4548 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4549  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4549 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4550  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4550 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4551  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4551 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4552  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4552 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4553  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4553 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4554  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4554 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4555  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4555 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4556  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4556 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4557  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4557 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4558  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4558 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4559  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4559 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4560  (.I0(\edb_top_inst/la0/GEN_PROBE[6].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[6].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4560 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4561  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4561 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4562  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4562 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4563  (.I0(\edb_top_inst/la0/GEN_PROBE[7].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4563 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4564  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4564 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4565  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3076 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4565 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4566  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3077 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4566 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4567  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4567 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4568  (.I0(\edb_top_inst/n3077 ), .I1(\edb_top_inst/n3076 ), 
            .I2(\edb_top_inst/n3078 ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4568 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4569  (.I0(\edb_top_inst/n2869 ), .I1(\edb_top_inst/n2870 ), 
            .O(\edb_top_inst/la0/n9630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4569 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4570  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4570 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4571  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4571 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4572  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), .O(\edb_top_inst/n3079 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4572 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4573  (.I0(\edb_top_inst/n3079 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), .O(\edb_top_inst/n3080 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4573 .LUTMASK = 16'h7171;
    EFX_LUT4 \edb_top_inst/LUT__4574  (.I0(\edb_top_inst/n3080 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), .O(\edb_top_inst/n3081 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4574 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4575  (.I0(\edb_top_inst/n3081 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), .O(\edb_top_inst/n3082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4575 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4576  (.I0(\edb_top_inst/n3082 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), .O(\edb_top_inst/n3083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4576 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4577  (.I0(\edb_top_inst/n3083 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), .O(\edb_top_inst/n3084 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4577 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4578  (.I0(\edb_top_inst/n3084 ), .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4578 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4579  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3085 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4579 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4580  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n3086 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4580 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4581  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3087 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4581 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4582  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3088 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4582 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4583  (.I0(\edb_top_inst/n3085 ), .I1(\edb_top_inst/n3086 ), 
            .I2(\edb_top_inst/n3087 ), .I3(\edb_top_inst/n3088 ), .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4583 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4584  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3089 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4584 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4585  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3090 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4585 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4586  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n3091 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4586 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4587  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3092 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4587 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4588  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3093 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4588 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4589  (.I0(\edb_top_inst/n3090 ), .I1(\edb_top_inst/n3091 ), 
            .I2(\edb_top_inst/n3092 ), .I3(\edb_top_inst/n3093 ), .O(\edb_top_inst/n3094 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4589 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4590  (.I0(\edb_top_inst/n3089 ), .I1(\edb_top_inst/n3094 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3095 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4590 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__4591  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3096 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4591 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4592  (.I0(\edb_top_inst/n3096 ), .I1(\edb_top_inst/n3095 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4592 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4593  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4593 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4594  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4594 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4595  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4595 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4596  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4596 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4597  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4597 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4598  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4598 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4599  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4599 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4600  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4600 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4601  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4601 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4602  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4602 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4603  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4603 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4604  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4604 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4605  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4605 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4606  (.I0(\edb_top_inst/la0/GEN_PROBE[8].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4606 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4607  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4607 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4608  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4608 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4609  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), .O(\edb_top_inst/n3097 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4609 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4610  (.I0(\edb_top_inst/n3097 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), .O(\edb_top_inst/n3098 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4610 .LUTMASK = 16'h7171;
    EFX_LUT4 \edb_top_inst/LUT__4611  (.I0(\edb_top_inst/n3098 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), .O(\edb_top_inst/n3099 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4611 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4612  (.I0(\edb_top_inst/n3099 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), .O(\edb_top_inst/n3100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4612 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4613  (.I0(\edb_top_inst/n3100 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), .O(\edb_top_inst/n3101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4613 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4614  (.I0(\edb_top_inst/n3101 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), .O(\edb_top_inst/n3102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4614 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4615  (.I0(\edb_top_inst/n3102 ), .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4615 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4616  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n3103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4616 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4617  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n3104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4617 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4618  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4618 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4619  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n3106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4619 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4620  (.I0(\edb_top_inst/n3103 ), .I1(\edb_top_inst/n3104 ), 
            .I2(\edb_top_inst/n3105 ), .I3(\edb_top_inst/n3106 ), .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4620 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4621  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n3107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4621 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4622  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n3108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4622 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4623  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n3109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4623 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4624  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n3110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4624 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4625  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n3111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4625 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4626  (.I0(\edb_top_inst/n3108 ), .I1(\edb_top_inst/n3109 ), 
            .I2(\edb_top_inst/n3110 ), .I3(\edb_top_inst/n3111 ), .O(\edb_top_inst/n3112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4626 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4627  (.I0(\edb_top_inst/n3107 ), .I1(\edb_top_inst/n3112 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4627 .LUTMASK = 16'h5c3f;
    EFX_LUT4 \edb_top_inst/LUT__4628  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n3114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4628 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4629  (.I0(\edb_top_inst/n3114 ), .I1(\edb_top_inst/n3113 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4629 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__4630  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4630 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4631  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4631 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4632  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4632 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4633  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4633 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4634  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4634 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4635  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4635 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4636  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4636 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4637  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4637 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4638  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4638 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4639  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4639 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4640  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4640 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4641  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4641 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4642  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4642 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4643  (.I0(\edb_top_inst/la0/GEN_PROBE[9].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4643 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4644  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4644 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4645  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4645 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4646  (.I0(\edb_top_inst/la0/GEN_PROBE[10].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4646 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4647  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4647 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4648  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4648 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4649  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4649 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4650  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4650 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4651  (.I0(\edb_top_inst/n3116 ), .I1(\edb_top_inst/n3115 ), 
            .I2(\edb_top_inst/n3117 ), .I3(\edb_top_inst/la0/GEN_PROBE[10].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4651 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4652  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4652 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4653  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4653 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4654  (.I0(\edb_top_inst/la0/GEN_PROBE[11].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4654 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4655  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4655 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4656  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n3118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4656 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4657  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4657 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__4658  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n3120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4658 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4659  (.I0(\edb_top_inst/n3119 ), .I1(\edb_top_inst/n3118 ), 
            .I2(\edb_top_inst/n3120 ), .I3(\edb_top_inst/la0/GEN_PROBE[11].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4659 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__4660  (.I0(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4660 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4661  (.I0(\edb_top_inst/la0/la_trig_mask[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4661 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4662  (.I0(\edb_top_inst/la0/la_trig_mask[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4662 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4663  (.I0(\edb_top_inst/la0/la_trig_mask[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[4] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4663 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4664  (.I0(\edb_top_inst/n3121 ), .I1(\edb_top_inst/n3122 ), 
            .I2(\edb_top_inst/n3123 ), .I3(\edb_top_inst/n3124 ), .O(\edb_top_inst/n3125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4664 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4665  (.I0(\edb_top_inst/la0/la_trig_mask[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4665 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4666  (.I0(\edb_top_inst/la0/la_trig_mask[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n3127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4666 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4667  (.I0(\edb_top_inst/n3125 ), .I1(\edb_top_inst/n3126 ), 
            .I2(\edb_top_inst/n3127 ), .O(\edb_top_inst/n3128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4667 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4668  (.I0(\edb_top_inst/la0/GEN_PROBE[11].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[11] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[4] ), .O(\edb_top_inst/n3129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4668 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4669  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[0] ), .O(\edb_top_inst/n3130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4669 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4670  (.I0(\edb_top_inst/la0/GEN_PROBE[5].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[5] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[3] ), .O(\edb_top_inst/n3131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4670 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4671  (.I0(\edb_top_inst/la0/GEN_PROBE[8].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[1] ), .O(\edb_top_inst/n3132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4671 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4672  (.I0(\edb_top_inst/n3129 ), .I1(\edb_top_inst/n3130 ), 
            .I2(\edb_top_inst/n3131 ), .I3(\edb_top_inst/n3132 ), .O(\edb_top_inst/n3133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4672 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4673  (.I0(\edb_top_inst/la0/GEN_PROBE[9].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[9] ), .O(\edb_top_inst/n3134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4673 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4674  (.I0(\edb_top_inst/la0/GEN_PROBE[10].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[10] ), .I2(\edb_top_inst/la0/GEN_PROBE[6].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[6] ), .O(\edb_top_inst/n3135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4674 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4675  (.I0(\edb_top_inst/la0/GEN_PROBE[7].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[7] ), .I2(\edb_top_inst/n3134 ), 
            .I3(\edb_top_inst/n3135 ), .O(\edb_top_inst/n3136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4675 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__4676  (.I0(\edb_top_inst/n3133 ), .I1(\edb_top_inst/n3136 ), 
            .I2(\edb_top_inst/n3128 ), .I3(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .O(\edb_top_inst/n3137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4676 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__4677  (.I0(\edb_top_inst/n3128 ), .I1(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .I2(\edb_top_inst/n3137 ), .O(\edb_top_inst/la0/trigger_tu/n89 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc1c1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4677 .LUTMASK = 16'hc1c1;
    EFX_LUT4 \edb_top_inst/LUT__4678  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .I2(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n3138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4678 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4679  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[6] ), 
            .O(\edb_top_inst/n3139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4679 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4680  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .I2(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[10] ), .O(\edb_top_inst/n3140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4680 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4681  (.I0(\edb_top_inst/n3138 ), .I1(\edb_top_inst/n3139 ), 
            .I2(\edb_top_inst/n3140 ), .O(\edb_top_inst/n3141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4681 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4682  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[14] ), .I2(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n3142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4682 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4683  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[12] ), .I2(\edb_top_inst/n3141 ), 
            .I3(\edb_top_inst/n3142 ), .O(\edb_top_inst/n3143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4683 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4684  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4684 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__4685  (.I0(\edb_top_inst/n3144 ), .I1(\edb_top_inst/n3143 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4685 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4686  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[10] ), .O(\edb_top_inst/n3146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4686 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4687  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .I2(\edb_top_inst/n3138 ), 
            .I3(\edb_top_inst/n3139 ), .O(\edb_top_inst/n3147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4687 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4688  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/n3146 ), .I2(\edb_top_inst/n3147 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .O(\edb_top_inst/n3148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4688 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4689  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/n3141 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[11] ), .O(\edb_top_inst/n3149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4689 .LUTMASK = 16'heb7e;
    EFX_LUT4 \edb_top_inst/LUT__4690  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n3150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4690 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4691  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n3151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4691 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4692  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/n3150 ), .I2(\edb_top_inst/n3151 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .O(\edb_top_inst/n3152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4692 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4693  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .O(\edb_top_inst/n3153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4693 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__4694  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n3154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4694 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4695  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/n3138 ), 
            .I3(\edb_top_inst/n3154 ), .O(\edb_top_inst/n3155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4695 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__4696  (.I0(\edb_top_inst/n3152 ), .I1(\edb_top_inst/n3153 ), 
            .I2(\edb_top_inst/n3155 ), .I3(\edb_top_inst/n3142 ), .O(\edb_top_inst/n3156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4696 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4697  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .O(\edb_top_inst/n3157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4697 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4698  (.I0(\edb_top_inst/n3138 ), .I1(\edb_top_inst/n3139 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[7] ), .I3(\edb_top_inst/n3157 ), 
            .O(\edb_top_inst/n3158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4698 .LUTMASK = 16'h8700;
    EFX_LUT4 \edb_top_inst/LUT__4699  (.I0(\edb_top_inst/n3138 ), .I1(\edb_top_inst/n3139 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[7] ), .I3(\edb_top_inst/n3157 ), 
            .O(\edb_top_inst/n3159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8ff7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4699 .LUTMASK = 16'h8ff7;
    EFX_LUT4 \edb_top_inst/LUT__4700  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n3160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4700 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4701  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/n3160 ), .I2(\edb_top_inst/n3138 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n3161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4701 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4702  (.I0(\edb_top_inst/n3159 ), .I1(\edb_top_inst/n3158 ), 
            .I2(\edb_top_inst/n3161 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .O(\edb_top_inst/n3162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4702 .LUTMASK = 16'h050c;
    EFX_LUT4 \edb_top_inst/LUT__4703  (.I0(\edb_top_inst/n3148 ), .I1(\edb_top_inst/n3149 ), 
            .I2(\edb_top_inst/n3156 ), .I3(\edb_top_inst/n3162 ), .O(\edb_top_inst/n3163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4703 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4704  (.I0(\edb_top_inst/n3163 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3145 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n3164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4704 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4705  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n3165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4705 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4706  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4706 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4707  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[8] ), 
            .O(\edb_top_inst/n3167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4707 .LUTMASK = 16'hf40b;
    EFX_LUT4 \edb_top_inst/LUT__4708  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4708 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4709  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4709 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4710  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/n3169 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[14] ), 
            .O(\edb_top_inst/n3170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf807, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4710 .LUTMASK = 16'hf807;
    EFX_LUT4 \edb_top_inst/LUT__4711  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4711 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4712  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4712 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4713  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/n3171 ), 
            .I2(\edb_top_inst/n3172 ), .O(\edb_top_inst/n3173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4713 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4714  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/la0/la_window_depth[4] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n3174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4714 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4715  (.I0(\edb_top_inst/n3174 ), .I1(\edb_top_inst/n3173 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[6] ), .I3(\edb_top_inst/n3170 ), 
            .O(\edb_top_inst/n3175 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4715 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__4716  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ffc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4716 .LUTMASK = 16'h6ffc;
    EFX_LUT4 \edb_top_inst/LUT__4717  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/n3176 ), 
            .I3(\edb_top_inst/n3171 ), .O(\edb_top_inst/n3177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4717 .LUTMASK = 16'hf077;
    EFX_LUT4 \edb_top_inst/LUT__4718  (.I0(\edb_top_inst/n3177 ), .I1(\edb_top_inst/n3175 ), 
            .I2(\edb_top_inst/n3167 ), .O(\edb_top_inst/n3178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4718 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4719  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/n3165 ), .O(\edb_top_inst/n3179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4719 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4720  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4720 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4721  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[13] ), .I2(\edb_top_inst/n3180 ), 
            .O(\edb_top_inst/n3181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4721 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4722  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n3182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4722 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4723  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n3171 ), .I3(\edb_top_inst/la0/la_trig_pos[4] ), 
            .O(\edb_top_inst/n3183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4723 .LUTMASK = 16'h4fb0;
    EFX_LUT4 \edb_top_inst/LUT__4724  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[13] ), .O(\edb_top_inst/n3184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f82, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4724 .LUTMASK = 16'h7f82;
    EFX_LUT4 \edb_top_inst/LUT__4725  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4725 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4726  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/n3184 ), .I3(\edb_top_inst/la0/la_trig_pos[9] ), 
            .O(\edb_top_inst/n3186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4726 .LUTMASK = 16'h0c0b;
    EFX_LUT4 \edb_top_inst/LUT__4727  (.I0(\edb_top_inst/n3186 ), .I1(\edb_top_inst/n3181 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n3183 ), 
            .O(\edb_top_inst/n3187 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4727 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4728  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/n3169 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[12] ), 
            .O(\edb_top_inst/n3188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bf4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4728 .LUTMASK = 16'h0bf4;
    EFX_LUT4 \edb_top_inst/LUT__4729  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n3172 ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[2] ), .O(\edb_top_inst/n3189 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4729 .LUTMASK = 16'h40bf;
    EFX_LUT4 \edb_top_inst/LUT__4730  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4730 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4731  (.I0(\edb_top_inst/n3189 ), .I1(\edb_top_inst/n3190 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n3191 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4731 .LUTMASK = 16'he7e7;
    EFX_LUT4 \edb_top_inst/LUT__4732  (.I0(\edb_top_inst/n3169 ), .I1(\edb_top_inst/la0/la_window_depth[4] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[15] ), .I3(\edb_top_inst/la0/la_trig_pos[11] ), 
            .O(\edb_top_inst/n3192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4732 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__4733  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[0] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4733 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__4734  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4734 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4735  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/n3194 ), 
            .I2(\edb_top_inst/n3171 ), .O(\edb_top_inst/n3195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4735 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4736  (.I0(\edb_top_inst/n3192 ), .I1(\edb_top_inst/n3193 ), 
            .I2(\edb_top_inst/n3195 ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n3196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4736 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__4737  (.I0(\edb_top_inst/n3188 ), .I1(\edb_top_inst/n3191 ), 
            .I2(\edb_top_inst/n3187 ), .I3(\edb_top_inst/n3196 ), .O(\edb_top_inst/n3197 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4737 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4738  (.I0(\edb_top_inst/n3165 ), .I1(\edb_top_inst/n3178 ), 
            .I2(\edb_top_inst/n3197 ), .I3(\edb_top_inst/n3179 ), .O(\edb_top_inst/n3198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4738 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4739  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3198 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/n3164 ), .O(\edb_top_inst/n3199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4739 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__4740  (.I0(\edb_top_inst/n3194 ), .I1(\edb_top_inst/n3168 ), 
            .O(\edb_top_inst/n3200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4740 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4741  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4741 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__4742  (.I0(\edb_top_inst/n3201 ), .I1(\edb_top_inst/n3166 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4742 .LUTMASK = 16'h0a03;
    EFX_LUT4 \edb_top_inst/LUT__4743  (.I0(\edb_top_inst/n3200 ), .I1(\edb_top_inst/n3202 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .O(\edb_top_inst/n3203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4743 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4744  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/n3168 ), 
            .O(\edb_top_inst/n3204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4744 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4745  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/n3172 ), 
            .O(\edb_top_inst/n3205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4745 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__4746  (.I0(\edb_top_inst/n3204 ), .I1(\edb_top_inst/n3205 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .O(\edb_top_inst/n3206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4746 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4747  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I3(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3207 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdcf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4747 .LUTMASK = 16'hbdcf;
    EFX_LUT4 \edb_top_inst/LUT__4748  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4748 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4749  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3209 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4749 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4750  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3209 ), 
            .O(\edb_top_inst/n3210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4750 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4751  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n3185 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4751 .LUTMASK = 16'h0c0b;
    EFX_LUT4 \edb_top_inst/LUT__4752  (.I0(\edb_top_inst/n3210 ), .I1(\edb_top_inst/n3211 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .O(\edb_top_inst/n3212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4752 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__4753  (.I0(\edb_top_inst/n3207 ), .I1(\edb_top_inst/n3208 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I3(\edb_top_inst/n3212 ), 
            .O(\edb_top_inst/n3213 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4753 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__4754  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n3166 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4754 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4755  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3182 ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n3215 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4551, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4755 .LUTMASK = 16'h4551;
    EFX_LUT4 \edb_top_inst/LUT__4756  (.I0(\edb_top_inst/n3214 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .I3(\edb_top_inst/n3215 ), 
            .O(\edb_top_inst/n3216 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4756 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__4757  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n3171 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n3217 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4757 .LUTMASK = 16'h4fb0;
    EFX_LUT4 \edb_top_inst/LUT__4758  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3173 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), .I3(\edb_top_inst/n3217 ), 
            .O(\edb_top_inst/n3218 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3edf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4758 .LUTMASK = 16'h3edf;
    EFX_LUT4 \edb_top_inst/LUT__4759  (.I0(\edb_top_inst/n3216 ), .I1(\edb_top_inst/n3218 ), 
            .O(\edb_top_inst/n3219 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4759 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4760  (.I0(\edb_top_inst/n3203 ), .I1(\edb_top_inst/n3206 ), 
            .I2(\edb_top_inst/n3213 ), .I3(\edb_top_inst/n3219 ), .O(\edb_top_inst/n3220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4760 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4761  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), .I3(\edb_top_inst/n3172 ), 
            .O(\edb_top_inst/n3221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4761 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__4762  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I3(\edb_top_inst/n3190 ), .O(\edb_top_inst/n3222 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4762 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__4763  (.I0(\edb_top_inst/n3221 ), .I1(\edb_top_inst/n3222 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .I3(\edb_top_inst/n3209 ), 
            .O(\edb_top_inst/n3223 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4763 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__4764  (.I0(\edb_top_inst/n3214 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .O(\edb_top_inst/n3224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4764 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4765  (.I0(\edb_top_inst/n3194 ), .I1(\edb_top_inst/n3171 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .O(\edb_top_inst/n3225 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4765 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4766  (.I0(\edb_top_inst/n3201 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .O(\edb_top_inst/n3226 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf40b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4766 .LUTMASK = 16'hf40b;
    EFX_LUT4 \edb_top_inst/LUT__4767  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n3171 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .O(\edb_top_inst/n3227 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4767 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__4768  (.I0(\edb_top_inst/n3225 ), .I1(\edb_top_inst/n3217 ), 
            .I2(\edb_top_inst/n3226 ), .I3(\edb_top_inst/n3227 ), .O(\edb_top_inst/n3228 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4768 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4769  (.I0(\edb_top_inst/n3169 ), .I1(\edb_top_inst/n3182 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n3229 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4769 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4770  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n3185 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n3230 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4770 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4771  (.I0(\edb_top_inst/n3229 ), .I1(\edb_top_inst/n3230 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .O(\edb_top_inst/n3231 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4771 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__4772  (.I0(\edb_top_inst/n3223 ), .I1(\edb_top_inst/n3224 ), 
            .I2(\edb_top_inst/n3228 ), .I3(\edb_top_inst/n3231 ), .O(\edb_top_inst/n3232 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4772 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4773  (.I0(\edb_top_inst/n3204 ), .I1(\edb_top_inst/n3205 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[3] ), .I3(\edb_top_inst/la0/la_trig_pos[2] ), 
            .O(\edb_top_inst/n3233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4773 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4774  (.I0(\edb_top_inst/n3200 ), .I1(\edb_top_inst/n3202 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[11] ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n3234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hedf3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4774 .LUTMASK = 16'hedf3;
    EFX_LUT4 \edb_top_inst/LUT__4775  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n3180 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[15] ), .O(\edb_top_inst/n3235 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4775 .LUTMASK = 16'h3ff4;
    EFX_LUT4 \edb_top_inst/LUT__4776  (.I0(\edb_top_inst/n3235 ), .I1(\edb_top_inst/n3230 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[9] ), .I3(\edb_top_inst/n3167 ), 
            .O(\edb_top_inst/n3236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4776 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__4777  (.I0(\edb_top_inst/n3233 ), .I1(\edb_top_inst/n3234 ), 
            .I2(\edb_top_inst/n3175 ), .I3(\edb_top_inst/n3236 ), .O(\edb_top_inst/n3237 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4777 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4778  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4778 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4779  (.I0(\edb_top_inst/n3238 ), .I1(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[4] ), .I3(\edb_top_inst/n3210 ), 
            .O(\edb_top_inst/n3239 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4779 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__4780  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[1] ), .I3(\edb_top_inst/n3208 ), 
            .O(\edb_top_inst/n3240 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4780 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__4781  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n3169 ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3241 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4781 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4782  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/n3241 ), .I2(\edb_top_inst/la0/la_trig_pos[13] ), 
            .O(\edb_top_inst/n3242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4782 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__4783  (.I0(\edb_top_inst/n3239 ), .I1(\edb_top_inst/n3240 ), 
            .I2(\edb_top_inst/n3188 ), .I3(\edb_top_inst/n3242 ), .O(\edb_top_inst/n3243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4783 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4784  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/n3237 ), 
            .I2(\edb_top_inst/n3243 ), .O(\edb_top_inst/n3244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4784 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4785  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/la0/la_num_trigger[6] ), 
            .O(\edb_top_inst/n3245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4785 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4786  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[3] ), .O(\edb_top_inst/n3246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4786 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4787  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .O(\edb_top_inst/n3247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4787 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4788  (.I0(\edb_top_inst/n3245 ), .I1(\edb_top_inst/n3246 ), 
            .I2(\edb_top_inst/n3247 ), .O(\edb_top_inst/n3248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4788 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4789  (.I0(\edb_top_inst/la0/la_num_trigger[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), .O(\edb_top_inst/n3249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4789 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4790  (.I0(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), .I2(\edb_top_inst/n3248 ), 
            .I3(\edb_top_inst/n3249 ), .O(\edb_top_inst/n3250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd6bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4790 .LUTMASK = 16'hd6bf;
    EFX_LUT4 \edb_top_inst/LUT__4791  (.I0(\edb_top_inst/n3249 ), .I1(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I2(\edb_top_inst/la0/la_num_trigger[11] ), .I3(\edb_top_inst/la0/la_num_trigger[12] ), 
            .O(\edb_top_inst/n3251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe45, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4791 .LUTMASK = 16'hfe45;
    EFX_LUT4 \edb_top_inst/LUT__4792  (.I0(\edb_top_inst/la0/la_num_trigger[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .O(\edb_top_inst/n3252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4792 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4793  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .O(\edb_top_inst/n3253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4793 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4794  (.I0(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I1(\edb_top_inst/n3252 ), .I2(\edb_top_inst/n3253 ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .O(\edb_top_inst/n3254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4794 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4795  (.I0(\edb_top_inst/n3251 ), .I1(\edb_top_inst/n3254 ), 
            .O(\edb_top_inst/n3255 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4795 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4796  (.I0(\edb_top_inst/n3246 ), .I1(\edb_top_inst/n3245 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .I3(\edb_top_inst/la0/la_num_trigger[7] ), 
            .O(\edb_top_inst/n3256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h87f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4796 .LUTMASK = 16'h87f8;
    EFX_LUT4 \edb_top_inst/LUT__4797  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), .O(\edb_top_inst/n3257 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4797 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4798  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[9] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .O(\edb_top_inst/n3258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4798 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__4799  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/n3245 ), .I2(\edb_top_inst/n3246 ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .O(\edb_top_inst/n3259 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4799 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4800  (.I0(\edb_top_inst/n3258 ), .I1(\edb_top_inst/n3259 ), 
            .I2(\edb_top_inst/n3256 ), .I3(\edb_top_inst/n3257 ), .O(\edb_top_inst/n3260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4800 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4801  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .O(\edb_top_inst/n3261 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4801 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__4802  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/n3261 ), .I2(\edb_top_inst/n3246 ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .O(\edb_top_inst/n3262 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4802 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__4803  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/n3246 ), 
            .I3(\edb_top_inst/la0/la_num_trigger[6] ), .O(\edb_top_inst/n3263 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4803 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__4804  (.I0(\edb_top_inst/la0/la_num_trigger[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .O(\edb_top_inst/n3264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4804 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4805  (.I0(\edb_top_inst/la0/la_num_trigger[13] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[14] ), .I2(\edb_top_inst/la0/la_num_trigger[15] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[16] ), .O(\edb_top_inst/n3265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4805 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4806  (.I0(\edb_top_inst/n3264 ), .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I2(\edb_top_inst/la0/la_num_trigger[0] ), .I3(\edb_top_inst/n3265 ), 
            .O(\edb_top_inst/n3266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4806 .LUTMASK = 16'h1800;
    EFX_LUT4 \edb_top_inst/LUT__4807  (.I0(\edb_top_inst/n3262 ), .I1(\edb_top_inst/n3263 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I3(\edb_top_inst/n3266 ), 
            .O(\edb_top_inst/n3267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4807 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__4808  (.I0(\edb_top_inst/n3250 ), .I1(\edb_top_inst/n3260 ), 
            .I2(\edb_top_inst/n3255 ), .I3(\edb_top_inst/n3267 ), .O(\edb_top_inst/n3268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4808 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4809  (.I0(\edb_top_inst/n3268 ), .I1(\edb_top_inst/n3143 ), 
            .O(\edb_top_inst/n3269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4809 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4810  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4810 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4811  (.I0(\edb_top_inst/n3244 ), .I1(\edb_top_inst/n3220 ), 
            .I2(\edb_top_inst/n3269 ), .I3(\edb_top_inst/n3270 ), .O(\edb_top_inst/n3271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4811 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4812  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n3165 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4812 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__4813  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n3273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4813 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4814  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n3232 ), .I2(\edb_top_inst/n3272 ), .I3(\edb_top_inst/n3273 ), 
            .O(\edb_top_inst/n3274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4814 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4815  (.I0(\edb_top_inst/n3163 ), .I1(\edb_top_inst/n3273 ), 
            .I2(\edb_top_inst/n3274 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n3275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4815 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4816  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n3271 ), .I2(\edb_top_inst/n3199 ), .I3(\edb_top_inst/n3275 ), 
            .O(\edb_top_inst/la0/la_biu_inst/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4816 .LUTMASK = 16'h10ff;
    EFX_LUT4 \edb_top_inst/LUT__4817  (.I0(\edb_top_inst/n2825 ), .I1(\edb_top_inst/n2818 ), 
            .I2(\edb_top_inst/la0/biu_ready ), .O(\edb_top_inst/la0/la_biu_inst/n382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4817 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4818  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/n1315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4818 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4819  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), 
            .I3(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4819 .LUTMASK = 16'h00be;
    EFX_LUT4 \edb_top_inst/LUT__4820  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(\edb_top_inst/ceg_net351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4820 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4821  (.I0(\edb_top_inst/n3165 ), .I1(\edb_top_inst/n3178 ), 
            .I2(\edb_top_inst/n3197 ), .O(\edb_top_inst/n3276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4821 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4822  (.I0(\edb_top_inst/n3268 ), .I1(\edb_top_inst/n3165 ), 
            .O(\edb_top_inst/n3277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4822 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4823  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4823 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4824  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/n3277 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I3(\edb_top_inst/n3278 ), 
            .O(\edb_top_inst/n3279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4824 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4825  (.I0(\edb_top_inst/n2903 ), .I1(\edb_top_inst/n3276 ), 
            .I2(\edb_top_inst/n3271 ), .I3(\edb_top_inst/n3279 ), .O(\edb_top_inst/la0/la_biu_inst/n1300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4825 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__4826  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/n17781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4826 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4827  (.I0(\edb_top_inst/n3244 ), .I1(\edb_top_inst/n3220 ), 
            .I2(\edb_top_inst/n3269 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n3280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4827 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__4828  (.I0(\edb_top_inst/n3179 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4828 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4829  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4829 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__4830  (.I0(\edb_top_inst/n3276 ), .I1(\edb_top_inst/n3277 ), 
            .I2(\edb_top_inst/n3281 ), .I3(\edb_top_inst/n3282 ), .O(\edb_top_inst/n3283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4830 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4831  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/n2904 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4831 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4832  (.I0(\edb_top_inst/n3165 ), .I1(\edb_top_inst/n3278 ), 
            .I2(\edb_top_inst/n3268 ), .O(\edb_top_inst/n3285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4832 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4833  (.I0(\edb_top_inst/n3285 ), .I1(\edb_top_inst/n3284 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n3286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4833 .LUTMASK = 16'h0a0c;
    EFX_LUT4 \edb_top_inst/LUT__4834  (.I0(\edb_top_inst/n3280 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3283 ), .I3(\edb_top_inst/n3286 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4834 .LUTMASK = 16'hff0b;
    EFX_LUT4 \edb_top_inst/LUT__4835  (.I0(\edb_top_inst/n3144 ), .I1(\edb_top_inst/n3143 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n3163 ), 
            .O(\edb_top_inst/n3287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4835 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4836  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/n3165 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n3288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4836 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__4837  (.I0(\edb_top_inst/n2904 ), .I1(\edb_top_inst/n3232 ), 
            .I2(\edb_top_inst/n3288 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n3289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4837 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4838  (.I0(\edb_top_inst/n3287 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I3(\edb_top_inst/n3289 ), 
            .O(\edb_top_inst/n3290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4838 .LUTMASK = 16'hf100;
    EFX_LUT4 \edb_top_inst/LUT__4839  (.I0(\edb_top_inst/n3179 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n3277 ), .I3(\edb_top_inst/n3276 ), .O(\edb_top_inst/n3291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4839 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__4840  (.I0(\edb_top_inst/n3143 ), .I1(\edb_top_inst/n3268 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n3292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4840 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4841  (.I0(\edb_top_inst/n3288 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4841 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4842  (.I0(\edb_top_inst/n3244 ), .I1(\edb_top_inst/n3220 ), 
            .I2(\edb_top_inst/n3292 ), .I3(\edb_top_inst/n3293 ), .O(\edb_top_inst/n3294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4842 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__4843  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n3163 ), .I2(\edb_top_inst/n3273 ), .O(\edb_top_inst/n3295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4843 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4844  (.I0(\edb_top_inst/n3294 ), .I1(\edb_top_inst/n3291 ), 
            .I2(\edb_top_inst/n3290 ), .I3(\edb_top_inst/n3295 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4844 .LUTMASK = 16'hfff2;
    EFX_LUT4 \edb_top_inst/LUT__4845  (.I0(\edb_top_inst/la0/la_biu_inst/n382 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), 
            .O(\edb_top_inst/ceg_net348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4845 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__4846  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4846 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4847  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n3165 ), .I2(\edb_top_inst/n2903 ), .O(\edb_top_inst/la0/la_biu_inst/n2053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4847 .LUTMASK = 16'hbfbf;
    EFX_LUT4 \edb_top_inst/LUT__4848  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4848 .LUTMASK = 16'h05fc;
    EFX_LUT4 \edb_top_inst/LUT__4849  (.I0(\edb_top_inst/la0/la_biu_inst/n2053 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n3296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4849 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4850  (.I0(\edb_top_inst/n3232 ), .I1(\edb_top_inst/n3296 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4850 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4851  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n3297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4851 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4852  (.I0(\edb_top_inst/n3297 ), .I1(\edb_top_inst/la0/la_resetn ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4852 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4853  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4853 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4854  (.I0(\edb_top_inst/n3296 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/ceg_net355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4854 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4855  (.I0(\edb_top_inst/n2909 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4855 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4856  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[15] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4856 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4857  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[16] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4857 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4858  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[17] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4858 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4859  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[18] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4859 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4860  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[19] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4860 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4861  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[20] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4861 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4862  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[21] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4862 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4863  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[22] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4863 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4864  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[23] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4864 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4865  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[24] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4865 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4866  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[25] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4866 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4867  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[26] ), .I2(\edb_top_inst/n2909 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4867 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4868  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .O(\edb_top_inst/n3298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4868 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4869  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/n3298 ), 
            .I2(\edb_top_inst/n3215 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4869 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__4870  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3299 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4870 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__4871  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/n3299 ), 
            .O(\edb_top_inst/n3300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4871 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4872  (.I0(\edb_top_inst/n3180 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I3(\edb_top_inst/n3300 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4872 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4873  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n3301 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4873 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4874  (.I0(\edb_top_inst/n3168 ), .I1(\edb_top_inst/n3301 ), 
            .I2(\edb_top_inst/n3229 ), .O(\edb_top_inst/n3302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4874 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4875  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3303 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4875 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4876  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/n3303 ), 
            .I3(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3304 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4876 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4877  (.I0(\edb_top_inst/n3304 ), .I1(\edb_top_inst/n3172 ), 
            .I2(\edb_top_inst/n3302 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4877 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4878  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3305 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4878 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4879  (.I0(\edb_top_inst/n3305 ), .I1(\edb_top_inst/n3303 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4879 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4880  (.I0(\edb_top_inst/n3306 ), .I1(\edb_top_inst/n3172 ), 
            .O(\edb_top_inst/n3307 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4880 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4881  (.I0(\edb_top_inst/n3301 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I3(\edb_top_inst/n3307 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4881 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4882  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3308 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b04, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4882 .LUTMASK = 16'h0b04;
    EFX_LUT4 \edb_top_inst/LUT__4883  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3309 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4883 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4884  (.I0(\edb_top_inst/n3309 ), .I1(\edb_top_inst/n3305 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4884 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4885  (.I0(\edb_top_inst/n3310 ), .I1(\edb_top_inst/n3298 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4885 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__4886  (.I0(\edb_top_inst/n3308 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I2(\edb_top_inst/n3311 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4886 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4887  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4887 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4888  (.I0(\edb_top_inst/n3312 ), .I1(\edb_top_inst/n3309 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4888 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4889  (.I0(\edb_top_inst/n3299 ), .I1(\edb_top_inst/n3313 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4889 .LUTMASK = 16'ha300;
    EFX_LUT4 \edb_top_inst/LUT__4890  (.I0(\edb_top_inst/n3238 ), .I1(\edb_top_inst/n3308 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I3(\edb_top_inst/n3314 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4890 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4891  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/n3308 ), .O(\edb_top_inst/n3315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4891 .LUTMASK = 16'hd700;
    EFX_LUT4 \edb_top_inst/LUT__4892  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4892 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4893  (.I0(\edb_top_inst/n3316 ), .I1(\edb_top_inst/n3312 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4893 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4894  (.I0(\edb_top_inst/n3317 ), .I1(\edb_top_inst/n3304 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4894 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4895  (.I0(\edb_top_inst/n3315 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I2(\edb_top_inst/n3318 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4895 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4896  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n3182 ), .I2(\edb_top_inst/n3308 ), .O(\edb_top_inst/n3319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4896 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4897  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4897 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4898  (.I0(\edb_top_inst/n3320 ), .I1(\edb_top_inst/n3316 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4898 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4899  (.I0(\edb_top_inst/n3321 ), .I1(\edb_top_inst/n3306 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4899 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4900  (.I0(\edb_top_inst/n3319 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I2(\edb_top_inst/n3322 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4900 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4901  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4901 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4902  (.I0(\edb_top_inst/n3323 ), .I1(\edb_top_inst/n3320 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4902 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4903  (.I0(\edb_top_inst/n3324 ), .I1(\edb_top_inst/n3298 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4903 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__4904  (.I0(\edb_top_inst/n3310 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n3325 ), 
            .O(\edb_top_inst/n3326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4904 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4905  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I3(\edb_top_inst/n3326 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4905 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4906  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4906 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4907  (.I0(\edb_top_inst/n3327 ), .I1(\edb_top_inst/n3323 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4907 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4908  (.I0(\edb_top_inst/n3328 ), .I1(\edb_top_inst/n3299 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n3329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4908 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__4909  (.I0(\edb_top_inst/n3313 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n3329 ), 
            .O(\edb_top_inst/n3330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4909 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__4910  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I3(\edb_top_inst/n3330 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4910 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4911  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4911 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4912  (.I0(\edb_top_inst/n3331 ), .I1(\edb_top_inst/n3327 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4912 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4913  (.I0(\edb_top_inst/n3332 ), .I1(\edb_top_inst/n3317 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4913 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4914  (.I0(\edb_top_inst/n3304 ), .I1(\edb_top_inst/n3194 ), 
            .I2(\edb_top_inst/la0/la_window_depth[3] ), .I3(\edb_top_inst/n3333 ), 
            .O(\edb_top_inst/n3334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4914 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4915  (.I0(\edb_top_inst/n3201 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I3(\edb_top_inst/n3334 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4915 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__4916  (.I0(\edb_top_inst/n3182 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n3335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4916 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4917  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n3336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4917 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4918  (.I0(\edb_top_inst/n3336 ), .I1(\edb_top_inst/n3331 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n3337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4918 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4919  (.I0(\edb_top_inst/n3337 ), .I1(\edb_top_inst/n3321 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n3171 ), 
            .O(\edb_top_inst/n3338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4919 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__4920  (.I0(\edb_top_inst/n3306 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/n3194 ), .I3(\edb_top_inst/n3338 ), .O(\edb_top_inst/n3339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4920 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__4921  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] ), 
            .I1(\edb_top_inst/n3308 ), .I2(\edb_top_inst/n3335 ), .I3(\edb_top_inst/n3339 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4921 .LUTMASK = 16'h80ff;
    EFX_LUT4 \edb_top_inst/LUT__4922  (.I0(\edb_top_inst/n3172 ), .I1(\edb_top_inst/n3298 ), 
            .I2(\edb_top_inst/n3215 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4922 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__4923  (.I0(\edb_top_inst/n3180 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I3(\edb_top_inst/n3300 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4923 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4924  (.I0(\edb_top_inst/n3304 ), .I1(\edb_top_inst/n3172 ), 
            .I2(\edb_top_inst/n3302 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4924 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4925  (.I0(\edb_top_inst/n3301 ), .I1(\edb_top_inst/n3229 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I3(\edb_top_inst/n3307 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4925 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4926  (.I0(\edb_top_inst/n3308 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I2(\edb_top_inst/n3311 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4926 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4927  (.I0(\edb_top_inst/n3238 ), .I1(\edb_top_inst/n3308 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I3(\edb_top_inst/n3314 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4927 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4928  (.I0(\edb_top_inst/n3315 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I2(\edb_top_inst/n3318 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4928 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4929  (.I0(\edb_top_inst/n3319 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I2(\edb_top_inst/n3322 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4929 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4930  (.I0(\edb_top_inst/n3166 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I3(\edb_top_inst/n3326 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4930 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4931  (.I0(\edb_top_inst/n3185 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I3(\edb_top_inst/n3330 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4931 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4932  (.I0(\edb_top_inst/n3201 ), .I1(\edb_top_inst/n3319 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I3(\edb_top_inst/n3334 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4932 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__4933  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] ), 
            .I1(\edb_top_inst/n3308 ), .I2(\edb_top_inst/n3335 ), .I3(\edb_top_inst/n3339 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4933 .LUTMASK = 16'h80ff;
    EFX_LUT4 \edb_top_inst/LUT__4934  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n3340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fb8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4934 .LUTMASK = 16'h0fb8;
    EFX_LUT4 \edb_top_inst/LUT__4935  (.I0(\edb_top_inst/n3340 ), .I1(jtag_inst2_SEL), 
            .I2(jtag_inst2_UPDATE), .I3(\edb_top_inst/edb_user_dr[81] ), 
            .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4935 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4936  (.I0(jtag_inst2_SEL), .I1(jtag_inst2_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4936 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4937  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[1] ), .O(\edb_top_inst/n2739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4937 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4945  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i4_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4945 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4946  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i5_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4946 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4947  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i8_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4947 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4948  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i9_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4948 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4949  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i10_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4949 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4950  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i11_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4950 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4951  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i12_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4951 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4952  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i13_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4952 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4953  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i14_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4953 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4954  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i15_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4954 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4955  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i16_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4955 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4956  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i17_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4956 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4957  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i18_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4957 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4958  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i19_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4958 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4959  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i20_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4959 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4960  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i21_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4960 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4961  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i22_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4961 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4962  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i23_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4962 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4963  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i25_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4963 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4964  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i26_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4964 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4965  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i27_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4965 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4966  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i28_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4966 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4967  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i29_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4967 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4968  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i30_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4968 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4969  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i31_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4969 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4970  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i32_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4970 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4971  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i33_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4971 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4972  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i34_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4972 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4973  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i35_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4973 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4974  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i36_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4974 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4975  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i37_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4975 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4976  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i38_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4976 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4977  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i39_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4977 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__4978  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/dff_57/i40_pre ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4978 .LUTMASK = 16'h5555;
    EFX_LUT4 \edb_top_inst/LUT__3984  (.I0(\edb_top_inst/la0/crc_data_out[21] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n2758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3984 .LUTMASK = 16'h9009;
    EFX_ADD \edb_top_inst/la0/add_91/i1  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/n1249 ), .CI(1'b0), .O(\edb_top_inst/n67 ), 
            .CO(\edb_top_inst/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i2  (.I0(\edb_top_inst/la0/bit_count[1] ), 
            .I1(\edb_top_inst/la0/bit_count[0] ), .CI(1'b0), .O(\edb_top_inst/n69 ), 
            .CO(\edb_top_inst/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .CI(1'b0), 
            .O(\edb_top_inst/n73 ), .CO(\edb_top_inst/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n693 ), .CO(\edb_top_inst/n694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n695 ), .CO(\edb_top_inst/n696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .CI(1'b0), 
            .CO(\edb_top_inst/n697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[0] ), .CI(1'b0), .CO(\edb_top_inst/n698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(1'b1), .CI(n8454), .O(\edb_top_inst/n710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4673)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_43/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(1'b1), .CI(n8455), .O(\edb_top_inst/n711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4659)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/sub_18/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13  (.I0(\edb_top_inst/la0/la_sample_cnt[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n714 ), .O(\edb_top_inst/n712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n716 ), .O(\edb_top_inst/n713 ), 
            .CO(\edb_top_inst/n714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n718 ), .O(\edb_top_inst/n715 ), 
            .CO(\edb_top_inst/n716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n720 ), .O(\edb_top_inst/n717 ), 
            .CO(\edb_top_inst/n718 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n722 ), .O(\edb_top_inst/n719 ), 
            .CO(\edb_top_inst/n720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n724 ), .O(\edb_top_inst/n721 ), 
            .CO(\edb_top_inst/n722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n726 ), .O(\edb_top_inst/n723 ), 
            .CO(\edb_top_inst/n724 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n728 ), .O(\edb_top_inst/n725 ), 
            .CO(\edb_top_inst/n726 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n730 ), .O(\edb_top_inst/n727 ), 
            .CO(\edb_top_inst/n728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n732 ), .O(\edb_top_inst/n729 ), 
            .CO(\edb_top_inst/n730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n698 ), .O(\edb_top_inst/n731 ), 
            .CO(\edb_top_inst/n732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4675)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n735 ), .O(\edb_top_inst/n733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n737 ), .O(\edb_top_inst/n734 ), 
            .CO(\edb_top_inst/n735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n739 ), .O(\edb_top_inst/n736 ), 
            .CO(\edb_top_inst/n737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n741 ), .O(\edb_top_inst/n738 ), 
            .CO(\edb_top_inst/n739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n743 ), .O(\edb_top_inst/n740 ), 
            .CO(\edb_top_inst/n741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n745 ), .O(\edb_top_inst/n742 ), 
            .CO(\edb_top_inst/n743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n747 ), .O(\edb_top_inst/n744 ), 
            .CO(\edb_top_inst/n745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n749 ), .O(\edb_top_inst/n746 ), 
            .CO(\edb_top_inst/n747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n751 ), .O(\edb_top_inst/n748 ), 
            .CO(\edb_top_inst/n749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n753 ), .O(\edb_top_inst/n750 ), 
            .CO(\edb_top_inst/n751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n697 ), .O(\edb_top_inst/n752 ), 
            .CO(\edb_top_inst/n753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4661)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n841 ), .O(\edb_top_inst/n838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n843 ), .O(\edb_top_inst/n840 ), 
            .CO(\edb_top_inst/n841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n845 ), .O(\edb_top_inst/n842 ), 
            .CO(\edb_top_inst/n843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n847 ), .O(\edb_top_inst/n844 ), 
            .CO(\edb_top_inst/n845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n849 ), .O(\edb_top_inst/n846 ), 
            .CO(\edb_top_inst/n847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n851 ), .O(\edb_top_inst/n848 ), 
            .CO(\edb_top_inst/n849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n853 ), .O(\edb_top_inst/n850 ), 
            .CO(\edb_top_inst/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n855 ), .O(\edb_top_inst/n852 ), 
            .CO(\edb_top_inst/n853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n857 ), .O(\edb_top_inst/n854 ), 
            .CO(\edb_top_inst/n855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n696 ), .O(\edb_top_inst/n856 ), 
            .CO(\edb_top_inst/n857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4654)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1009 ), .O(\edb_top_inst/n1005 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1012 ), .O(\edb_top_inst/n1008 ), 
            .CO(\edb_top_inst/n1009 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1014 ), .O(\edb_top_inst/n1011 ), 
            .CO(\edb_top_inst/n1012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1016 ), .O(\edb_top_inst/n1013 ), 
            .CO(\edb_top_inst/n1014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1018 ), .O(\edb_top_inst/n1015 ), 
            .CO(\edb_top_inst/n1016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1020 ), .O(\edb_top_inst/n1017 ), 
            .CO(\edb_top_inst/n1018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1022 ), .O(\edb_top_inst/n1019 ), 
            .CO(\edb_top_inst/n1020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1024 ), .O(\edb_top_inst/n1021 ), 
            .CO(\edb_top_inst/n1022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1026 ), .O(\edb_top_inst/n1023 ), 
            .CO(\edb_top_inst/n1024 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n694 ), .O(\edb_top_inst/n1025 ), 
            .CO(\edb_top_inst/n1026 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4650)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1029 ), .O(\edb_top_inst/n1027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1031 ), .O(\edb_top_inst/n1028 ), 
            .CO(\edb_top_inst/n1029 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1033 ), .O(\edb_top_inst/n1030 ), 
            .CO(\edb_top_inst/n1031 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1035 ), .O(\edb_top_inst/n1032 ), 
            .CO(\edb_top_inst/n1033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1037 ), .O(\edb_top_inst/n1034 ), 
            .CO(\edb_top_inst/n1035 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1039 ), .O(\edb_top_inst/n1036 ), 
            .CO(\edb_top_inst/n1037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1041 ), .O(\edb_top_inst/n1038 ), 
            .CO(\edb_top_inst/n1039 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1043 ), .O(\edb_top_inst/n1040 ), 
            .CO(\edb_top_inst/n1041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1045 ), .O(\edb_top_inst/n1042 ), 
            .CO(\edb_top_inst/n1043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n74 ), .O(\edb_top_inst/n1044 ), 
            .CO(\edb_top_inst/n1045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i6  (.I0(\edb_top_inst/la0/bit_count[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1048 ), .O(\edb_top_inst/n1046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i5  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1050 ), .O(\edb_top_inst/n1047 ), 
            .CO(\edb_top_inst/n1048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i4  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1052 ), .O(\edb_top_inst/n1049 ), 
            .CO(\edb_top_inst/n1050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i3  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n70 ), .O(\edb_top_inst/n1051 ), 
            .CO(\edb_top_inst/n1052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3721)
    defparam \edb_top_inst/la0/add_100/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i27  (.I0(\edb_top_inst/la0/address_counter[26] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1065 ), .O(\edb_top_inst/n1062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i27 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i26  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1067 ), .O(\edb_top_inst/n1064 ), 
            .CO(\edb_top_inst/n1065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i26 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i25  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1069 ), .O(\edb_top_inst/n1066 ), 
            .CO(\edb_top_inst/n1067 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i24  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1071 ), .O(\edb_top_inst/n1068 ), 
            .CO(\edb_top_inst/n1069 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i23  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1073 ), .O(\edb_top_inst/n1070 ), 
            .CO(\edb_top_inst/n1071 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i22  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1075 ), .O(\edb_top_inst/n1072 ), 
            .CO(\edb_top_inst/n1073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i21  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1077 ), .O(\edb_top_inst/n1074 ), 
            .CO(\edb_top_inst/n1075 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i20  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1079 ), .O(\edb_top_inst/n1076 ), 
            .CO(\edb_top_inst/n1077 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i19  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1081 ), .O(\edb_top_inst/n1078 ), 
            .CO(\edb_top_inst/n1079 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i18  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1083 ), .O(\edb_top_inst/n1080 ), 
            .CO(\edb_top_inst/n1081 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i17  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1085 ), .O(\edb_top_inst/n1082 ), 
            .CO(\edb_top_inst/n1083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i16  (.I0(\edb_top_inst/la0/address_counter[15] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1087 ), .O(\edb_top_inst/n1084 ), 
            .CO(\edb_top_inst/n1085 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i15  (.I0(\edb_top_inst/la0/address_counter[14] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1089 ), .O(\edb_top_inst/n1086 ), 
            .CO(\edb_top_inst/n1087 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i14  (.I0(\edb_top_inst/la0/address_counter[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1091 ), .O(\edb_top_inst/n1088 ), 
            .CO(\edb_top_inst/n1089 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i13  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1093 ), .O(\edb_top_inst/n1090 ), 
            .CO(\edb_top_inst/n1091 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i12  (.I0(\edb_top_inst/la0/address_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1095 ), .O(\edb_top_inst/n1092 ), 
            .CO(\edb_top_inst/n1093 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i11  (.I0(\edb_top_inst/la0/address_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1097 ), .O(\edb_top_inst/n1094 ), 
            .CO(\edb_top_inst/n1095 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i10  (.I0(\edb_top_inst/la0/address_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1099 ), .O(\edb_top_inst/n1096 ), 
            .CO(\edb_top_inst/n1097 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i9  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1101 ), .O(\edb_top_inst/n1098 ), 
            .CO(\edb_top_inst/n1099 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i8  (.I0(\edb_top_inst/la0/address_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1103 ), .O(\edb_top_inst/n1100 ), 
            .CO(\edb_top_inst/n1101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i7  (.I0(\edb_top_inst/la0/address_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1105 ), .O(\edb_top_inst/n1102 ), 
            .CO(\edb_top_inst/n1103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i6  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1107 ), .O(\edb_top_inst/n1104 ), 
            .CO(\edb_top_inst/n1105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i5  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1109 ), .O(\edb_top_inst/n1106 ), 
            .CO(\edb_top_inst/n1107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i4  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/n2733 ), .CI(\edb_top_inst/n1111 ), .O(\edb_top_inst/n1108 ), 
            .CO(\edb_top_inst/n1109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i3  (.I0(\edb_top_inst/la0/address_counter[2] ), 
            .I1(\edb_top_inst/n2736 ), .CI(\edb_top_inst/n1113 ), .O(\edb_top_inst/n1110 ), 
            .CO(\edb_top_inst/n1111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i2  (.I0(\edb_top_inst/la0/address_counter[1] ), 
            .I1(\edb_top_inst/n2739 ), .CI(\edb_top_inst/n68 ), .O(\edb_top_inst/n1112 ), 
            .CO(\edb_top_inst/n1113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3694)
    defparam \edb_top_inst/la0/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i12  (.I0(\edb_top_inst/la0/address_counter[26] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1126 ), .O(\edb_top_inst/n1123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i11  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1128 ), .O(\edb_top_inst/n1125 ), 
            .CO(\edb_top_inst/n1126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i10  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1130 ), .O(\edb_top_inst/n1127 ), 
            .CO(\edb_top_inst/n1128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i9  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1132 ), .O(\edb_top_inst/n1129 ), 
            .CO(\edb_top_inst/n1130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i8  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1134 ), .O(\edb_top_inst/n1131 ), 
            .CO(\edb_top_inst/n1132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i7  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1136 ), .O(\edb_top_inst/n1133 ), 
            .CO(\edb_top_inst/n1134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i6  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1138 ), .O(\edb_top_inst/n1135 ), 
            .CO(\edb_top_inst/n1136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i5  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1143 ), .O(\edb_top_inst/n1137 ), 
            .CO(\edb_top_inst/n1138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i4  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1145 ), .O(\edb_top_inst/n1142 ), 
            .CO(\edb_top_inst/n1143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i3  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1147 ), .O(\edb_top_inst/n1144 ), 
            .CO(\edb_top_inst/n1145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i2  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(\edb_top_inst/la0/address_counter[15] ), .CI(1'b0), .O(\edb_top_inst/n1146 ), 
            .CO(\edb_top_inst/n1147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // D:/workspace/Efinix/Titanium/Ti180MIPI25GRxHDMIV101/work_dbg/debug_top.v(3693)
    defparam \edb_top_inst/la0/add_90/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i2 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__11266 (.I0(\MCsiRxController/MCsi2Decoder/wFtiRd[16] ), 
            .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), .I2(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .O(\MCsiRxController/MCsi2Decoder/n631 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h03e0 */ ;
    defparam LUT__11266.LUTMASK = 16'h03e0;
    EFX_LUT4 LUT__11267 (.I0(rSRST), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .O(\MCsiRxController/MCsi2Decoder/n633 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11267.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11268 (.I0(oTestPort[24]), .I1(oTestPort[0]), .O(\MCsiRxController/MCsi2Decoder/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11268.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11269 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[1] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .O(n8177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11269.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11270 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[4] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .O(n8178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11270.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11271 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[6] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .O(n8179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11271.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11272 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[8] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[9] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .O(n8180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11272.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11273 (.I0(n8177), .I1(n8178), .I2(n8179), .I3(n8180), 
            .O(n8181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11273.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11274 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[2] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rORP[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .O(n8182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11274.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11275 (.I0(n8181), .I1(n8182), .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRVd )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__11275.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__11276 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .O(n8183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11276.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11277 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .O(n8184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11277.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11278 (.I0(n8184), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(n8185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11278.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11279 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(n8183), .I2(n8185), .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(n8186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__11279.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__11280 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .O(n8187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11280.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11281 (.I0(n8185), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I3(n8187), .O(n8188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__11281.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__11282 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(n8189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11282.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11283 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(n8190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__11283.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__11284 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n8191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11284.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11285 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I2(n8191), .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(n8192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f */ ;
    defparam LUT__11285.LUTMASK = 16'hed3f;
    EFX_LUT4 LUT__11286 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n8193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11286.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11287 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .O(n8194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he33c */ ;
    defparam LUT__11287.LUTMASK = 16'he33c;
    EFX_LUT4 LUT__11288 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .O(n8195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11288.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11289 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(n8193), .I2(n8194), .I3(n8195), .O(n8196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__11289.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__11290 (.I0(n8192), .I1(n8196), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .O(n8197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001 */ ;
    defparam LUT__11290.LUTMASK = 16'h1001;
    EFX_LUT4 LUT__11291 (.I0(n8190), .I1(n8189), .I2(n8184), .I3(n8197), 
            .O(n8198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__11291.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__11292 (.I0(n8184), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(n8199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11292.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11293 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I1(n8183), .I2(n8199), .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(n8200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__11293.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__11294 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .O(n8201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11294.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11295 (.I0(n8191), .I1(n8201), .O(n8202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11295.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11296 (.I0(n8192), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(n8202), .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .O(n8203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__11296.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__11297 (.I0(n8199), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I3(n8187), .O(n8204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__11297.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__11298 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(n8205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__11298.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__11299 (.I0(n8205), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(n8193), .I3(n8195), .O(n8206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc8bf */ ;
    defparam LUT__11299.LUTMASK = 16'hc8bf;
    EFX_LUT4 LUT__11300 (.I0(n8184), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .O(n8207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11300.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11301 (.I0(n8190), .I1(n8189), .I2(n8206), .I3(n8207), 
            .O(n8208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__11301.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__11302 (.I0(n8200), .I1(n8203), .I2(n8204), .I3(n8208), 
            .O(n8209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11302.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11303 (.I0(n8188), .I1(n8186), .I2(n8198), .I3(n8209), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qFullAllmost )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__11303.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__11304 (.I0(\wHsDatatype[2] ), .I1(\wHsDatatype[3] ), .I2(\wHsDatatype[4] ), 
            .I3(\wHsDatatype[5] ), .O(n8210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__11304.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__11305 (.I0(n8210), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I3(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .O(n8211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff3 */ ;
    defparam LUT__11305.LUTMASK = 16'heff3;
    EFX_LUT4 LUT__11306 (.I0(n8211), .I1(rSRST), .I2(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .O(\MCsiRxController/MCsi2Decoder/n585 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__11306.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__11307 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .I3(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .O(\MCsiRxController/MCsi2Decoder/n604 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800 */ ;
    defparam LUT__11307.LUTMASK = 16'h1800;
    EFX_LUT4 LUT__11308 (.I0(\wHsWordCnt[11] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), 
            .I2(\wHsWordCnt[12] ), .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .O(n8212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11308.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11309 (.I0(\wHsWordCnt[11] ), .I1(\wHsWordCnt[12] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[11] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[10] ), .O(n8213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__11309.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__11310 (.I0(\wHsWordCnt[10] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[9] ), 
            .O(n8214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11310.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11311 (.I0(\wHsWordCnt[1] ), .I1(\wHsWordCnt[2] ), .I2(\wHsWordCnt[3] ), 
            .I3(\wHsWordCnt[4] ), .O(n8215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11311.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11312 (.I0(\wHsWordCnt[5] ), .I1(\wHsWordCnt[6] ), .I2(\wHsWordCnt[7] ), 
            .I3(\wHsWordCnt[8] ), .O(n8216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11312.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11313 (.I0(n8215), .I1(n8216), .O(n8217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11313.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11314 (.I0(\wHsWordCnt[9] ), .I1(n8214), .I2(n8217), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[8] ), .O(n8218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__11314.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__11315 (.I0(\wHsWordCnt[9] ), .I1(\wHsWordCnt[10] ), .I2(n8215), 
            .I3(n8216), .O(n8219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11315.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11316 (.I0(n8213), .I1(n8212), .I2(n8218), .I3(n8219), 
            .O(n8220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__11316.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__11317 (.I0(\wHsWordCnt[8] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[7] ), 
            .O(n8221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11317.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11318 (.I0(\wHsWordCnt[5] ), .I1(\wHsWordCnt[6] ), .I2(n8215), 
            .O(n8222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11318.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11319 (.I0(\wHsWordCnt[7] ), .I1(n8221), .I2(n8222), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[6] ), .O(n8223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__11319.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__11320 (.I0(\wHsWordCnt[6] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[5] ), 
            .O(n8224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11320.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11321 (.I0(n8224), .I1(n8215), .I2(\wHsWordCnt[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[4] ), .O(n8225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__11321.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__11322 (.I0(\wHsWordCnt[4] ), .I1(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[3] ), 
            .O(n8226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11322.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11323 (.I0(\wHsWordCnt[1] ), .I1(\wHsWordCnt[2] ), .O(n8227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11323.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11324 (.I0(\wHsWordCnt[3] ), .I1(n8226), .I2(n8227), 
            .I3(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[2] ), .O(n8228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__11324.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__11325 (.I0(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[0] ), 
            .I1(\wHsWordCnt[2] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[1] ), 
            .I3(\wHsWordCnt[1] ), .O(n8229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7 */ ;
    defparam LUT__11325.LUTMASK = 16'hbed7;
    EFX_LUT4 LUT__11326 (.I0(n8229), .I1(\wHsWordCnt[15] ), .I2(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .O(n8230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11326.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11327 (.I0(n8223), .I1(n8225), .I2(n8228), .I3(n8230), 
            .O(n8231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11327.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11328 (.I0(\wHsWordCnt[14] ), .I1(\wHsWordCnt[13] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] ), 
            .O(n8232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__11328.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__11329 (.I0(\wHsWordCnt[13] ), .I1(\wHsWordCnt[14] ), .I2(\MCsiRxController/MCsi2Decoder/rFrameWidthCnt[12] ), 
            .O(n8233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdbd */ ;
    defparam LUT__11329.LUTMASK = 16'hbdbd;
    EFX_LUT4 LUT__11330 (.I0(\wHsWordCnt[11] ), .I1(\wHsWordCnt[12] ), .I2(n8219), 
            .O(n8234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11330.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11331 (.I0(n8233), .I1(n8232), .I2(n8234), .O(n8235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__11331.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__11332 (.I0(n8235), .I1(n8231), .I2(n8220), .I3(rSRST), 
            .O(\MCsiRxController/MCsi2Decoder/qLineCntRst )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;
    defparam LUT__11332.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__11333 (.I0(n8183), .I1(n8187), .I2(n8195), .O(n8236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11333.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11334 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(n8237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11334.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11335 (.I0(n8202), .I1(n8236), .I2(n8189), .I3(n8237), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__11335.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__11336 (.I0(\MCsiRxController/MCsi2Decoder/wFtiEmp[0] ), 
            .I1(wCdcFifoFull), .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/equal_38/n19 ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11336.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11337 (.I0(n8233), .I1(n8232), .I2(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .I3(n8234), .O(n8238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h050c */ ;
    defparam LUT__11337.LUTMASK = 16'h050c;
    EFX_LUT4 LUT__11338 (.I0(n8238), .I1(n8220), .I2(n8231), .I3(n8211), 
            .O(\MCsiRxController/MCsi2Decoder/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__11338.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__11339 (.I0(\MCsiRxController/MCsi2Decoder/wFtiRvd[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), .I2(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), 
            .O(\MCsiRxController/MCsi2Decoder/n607 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c2c */ ;
    defparam LUT__11339.LUTMASK = 16'h2c2c;
    EFX_LUT4 LUT__11340 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11340.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11341 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11341.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11342 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11342.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11343 (.I0(n8193), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11343.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11344 (.I0(n8207), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11344.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11345 (.I0(n8207), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11345.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11346 (.I0(n8199), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n263 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11346.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11347 (.I0(n8199), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11347.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11348 (.I0(n8199), .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .O(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/n273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11348.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11349 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[8] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[8] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[9] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[9] ), 
            .O(n8239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11349.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11350 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[0] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rWA[0] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[1] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[1] ), 
            .O(n8240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11350.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11351 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[6] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[6] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[7] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[7] ), 
            .O(n8241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11351.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11352 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[4] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[4] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[5] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[5] ), 
            .O(n8242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11352.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11353 (.I0(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[2] ), 
            .I1(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/rRA[3] ), 
            .I3(\MCsiRxController/MCsi2Decoder/genblk1[0].Csi2DecoderDualClkFifo/rWA[3] ), 
            .O(n8243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11353.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11354 (.I0(n8240), .I1(n8241), .I2(n8242), .I3(n8243), 
            .O(n8244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11354.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11355 (.I0(n8244), .I1(n8239), .I2(\MCsiRxController/MCsi2Decoder/wFtiEmp[0] ), 
            .I3(wCdcFifoFull), .O(\MCsiRxController/MCsi2Decoder/genblk1[1].Csi2DecoderDualClkFifo/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__11355.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__11356 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .O(\MCsiRxController/MCsi2Decoder/equal_63/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__11356.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__11357 (.I0(\MCsiRxController/MCsi2Decoder/rHsSt[0] ), .I1(\MCsiRxController/MCsi2Decoder/rHsSt[2] ), 
            .I2(\MCsiRxController/MCsi2Decoder/rHsSt[1] ), .O(\MCsiRxController/MCsi2Decoder/equal_60/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__11357.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__11358 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] ), .O(n8245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11358.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11359 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .O(n8246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11359.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11360 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), .O(n8247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11360.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11361 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), .O(n8248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11361.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11362 (.I0(n8245), .I1(n8246), .I2(n8247), .I3(n8248), 
            .O(n8249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11362.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11363 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), .O(n8250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11363.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11364 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), .I2(n8249), 
            .I3(n8250), .O(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6fff */ ;
    defparam LUT__11364.LUTMASK = 16'h6fff;
    EFX_LUT4 LUT__11365 (.I0(\MCsiRxController/wFtiEmp[0] ), .I1(wVideofull), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/equal_75/n17 ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11365.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11366 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .O(n8251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11366.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11367 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I1(n8245), .I2(n8251), .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .O(n8252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__11367.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__11368 (.I0(n8246), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), .O(n8253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__11368.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__11369 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), 
            .O(n8254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11369.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11370 (.I0(n8254), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), .O(n8255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__11370.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__11371 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .I2(n8253), 
            .I3(n8255), .O(n8256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__11371.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__11372 (.I0(n8252), .I1(n8256), .O(n8257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11372.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11373 (.I0(n8251), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), 
            .O(n8258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11373.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11374 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I1(n8245), .I2(n8258), .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .O(n8259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__11374.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__11375 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(n8260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__11375.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__11376 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), .I2(n8246), 
            .O(n8261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787 */ ;
    defparam LUT__11376.LUTMASK = 16'h8787;
    EFX_LUT4 LUT__11377 (.I0(n8259), .I1(n8260), .I2(n8261), .I3(n8255), 
            .O(n8262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11377.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11378 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), .O(n8263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__11378.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__11379 (.I0(n8263), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), .O(n8264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__11379.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__11380 (.I0(n8257), .I1(n8249), .I2(n8262), .I3(n8264), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/qFullAllmost )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__11380.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__11381 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[3] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[3] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[6] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[6] ), .O(n8265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11381.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11382 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[4] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[4] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[7] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[7] ), .O(n8266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11382.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11383 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[0] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[2] ), .O(n8267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11383.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11384 (.I0(n8265), .I1(n8266), .I2(n8267), .O(n8268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11384.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11385 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[1] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[8] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[8] ), .O(n8269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11385.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11386 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rRA[5] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rORP[5] ), .I2(n8268), 
            .I3(n8269), .O(\MCsiRxController/genblk1[0].mVideoFIFO/qRVD )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6fff */ ;
    defparam LUT__11386.LUTMASK = 16'h6fff;
    EFX_LUT4 LUT__11387 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11387.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11388 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11388.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11389 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11389.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11390 (.I0(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[0] ), 
            .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[1] ), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[2] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[3] ), .O(n8270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11390.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11391 (.I0(n8270), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11391.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11392 (.I0(n8270), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11392.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11393 (.I0(n8270), .I1(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[4] ), 
            .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[5] ), .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[6] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11393.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11394 (.I0(n8251), .I1(n8270), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .O(\MCsiRxController/genblk1[0].mVideoFIFO/n466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11394.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11395 (.I0(n8251), .I1(n8270), .I2(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[7] ), 
            .I3(\MCsiRxController/genblk1[0].mVideoFIFO/rWA[8] ), .O(\MCsiRxController/genblk1[0].mVideoFIFO/n471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11395.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11396 (.I0(oTestPort[24]), .I1(n3048), .O(\MCsiRxController/n280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11396.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11397 (.I0(oTestPort[24]), .I1(n3046), .O(\MCsiRxController/n279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11397.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11398 (.I0(oTestPort[24]), .I1(n3044), .O(\MCsiRxController/n278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11398.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11399 (.I0(oTestPort[24]), .I1(n3042), .O(\MCsiRxController/n277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11399.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11400 (.I0(oTestPort[24]), .I1(n3040), .O(\MCsiRxController/n276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11400.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11401 (.I0(oTestPort[24]), .I1(n3038), .O(\MCsiRxController/n275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11401.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11402 (.I0(oTestPort[24]), .I1(n3036), .O(\MCsiRxController/n274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11402.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11403 (.I0(oTestPort[24]), .I1(n3034), .O(\MCsiRxController/n273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11403.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11404 (.I0(oTestPort[24]), .I1(n3032), .O(\MCsiRxController/n272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11404.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11405 (.I0(oTestPort[24]), .I1(n3030), .O(\MCsiRxController/n271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11405.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11406 (.I0(oTestPort[24]), .I1(n3028), .O(\MCsiRxController/n270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11406.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11407 (.I0(oTestPort[24]), .I1(n3026), .O(\MCsiRxController/n269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11407.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11408 (.I0(oTestPort[24]), .I1(n3024), .O(\MCsiRxController/n268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11408.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11409 (.I0(oTestPort[24]), .I1(n3022), .O(\MCsiRxController/n267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11409.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11410 (.I0(oTestPort[24]), .I1(n3021), .O(\MCsiRxController/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11410.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11411 (.I0(wVideoVd), .I1(\MVideoPostProcess/rVtgRstSel ), 
            .O(\MVideoPostProcess/qVtgRstCntCke )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11411.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11412 (.I0(\MVideoPostProcess/rVtgRstCnt[0] ), .I1(\MVideoPostProcess/rVtgRstCnt[1] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[2] ), .I3(\MVideoPostProcess/rVtgRstCnt[4] ), 
            .O(n8271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11412.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11413 (.I0(\MVideoPostProcess/rVtgRstCnt[3] ), .I1(\MVideoPostProcess/rVtgRstCnt[5] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[6] ), .I3(\MVideoPostProcess/rVtgRstCnt[10] ), 
            .O(n8272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11413.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11414 (.I0(\MVideoPostProcess/rVtgRstCnt[7] ), .I1(\MVideoPostProcess/rVtgRstCnt[8] ), 
            .I2(\MVideoPostProcess/rVtgRstCnt[9] ), .O(n8273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11414.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11415 (.I0(n8271), .I1(n8272), .I2(n8273), .O(\MVideoPostProcess/equal_18/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f7f */ ;
    defparam LUT__11415.LUTMASK = 16'h7f7f;
    EFX_LUT4 LUT__11416 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\~n1835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11416.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11417 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), 
            .O(n8274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11417.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11418 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), .O(n8275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11418.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11419 (.I0(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] ), 
            .I1(n8274), .I2(n8275), .O(n8276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11419.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11420 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_ack ), .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(n8277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11420.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11421 (.I0(n8276), .I1(n8277), .O(n8278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11421.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11422 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .I1(pll_inst1_LOCKED), .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I3(rBRST), .O(n8279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__11422.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__11423 (.I0(n8278), .I1(n8279), .O(ceg_net939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11423.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11424 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(n8276), .I2(n8277), .O(\MVideoPostProcess/inst_adv7511_config/n816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f1f */ ;
    defparam LUT__11424.LUTMASK = 16'h1f1f;
    EFX_LUT4 LUT__11425 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] ), .O(n8280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11425.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11426 (.I0(n8280), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] ), 
            .O(n8281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11426.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11427 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
            .I1(n8281), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] ), .O(n8282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11427.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11428 (.I0(n8282), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .I3(n8279), .O(\~ceg_net512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__11428.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__11429 (.I0(n8278), .I1(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11429.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11430 (.I0(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11430.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11431 (.I0(\MVideoPostProcess/inst_adv7511_config/n833 ), 
            .I1(n8279), .O(ceg_net995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11431.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11432 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11432.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11433 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_2P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/n1107 ), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_3P ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11433.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11434 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11434.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11435 (.I0(rBRST), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(ceg_net479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11435.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11436 (.I0(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(ceg_net43)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11436.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11437 (.I0(ceg_net479), .I1(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(n8283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11437.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11438 (.I0(\MVideoPostProcess/inst_adv7511_config/w_ack ), 
            .I1(n8276), .I2(n8283), .I3(\~ceg_net512 ), .O(ceg_net1327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__11438.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__11439 (.I0(rBRST), .I1(\MVideoPostProcess/inst_adv7511_config/n1107 ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n1243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11439.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11440 (.I0(iAdv7511Scl), .I1(oAdv7511SclOe), .I2(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .O(n8284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__11440.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__11441 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .O(n8285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11441.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11442 (.I0(n8285), .I1(n8284), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n8286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__11442.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__11443 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n8287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11443.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11444 (.I0(n8286), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(n8287), .O(n8288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__11444.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__11445 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(n8288), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11445.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11446 (.I0(n8287), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n8289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11446.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11447 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(n8289), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11447.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11448 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(n8287), .O(n8290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff0 */ ;
    defparam LUT__11448.LUTMASK = 16'heff0;
    EFX_LUT4 LUT__11449 (.I0(n8290), .I1(n8285), .I2(n8287), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(ceg_net1087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__11449.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__11450 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I2(oAdv7511SdaOe), .O(n8291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__11450.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__11451 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .I1(iAdv7511Sda), .I2(n8285), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n8292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__11451.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__11452 (.I0(n8292), .I1(n8291), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n8293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11452.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11453 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] ), 
            .O(n8294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11453.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11454 (.I0(n8285), .I1(n8294), .O(n8295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11454.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11455 (.I0(\MVideoPostProcess/inst_adv7511_config/r_last_1P ), 
            .I1(oAdv7511SdaOe), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(n8295), .O(n8296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a03 */ ;
    defparam LUT__11455.LUTMASK = 16'h0a03;
    EFX_LUT4 LUT__11456 (.I0(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n8297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__11456.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__11457 (.I0(n8285), .I1(n8297), .I2(n8291), .O(n8298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__11457.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__11458 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n8299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11458.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11459 (.I0(n8296), .I1(n8298), .I2(n8299), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n8300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11459.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11460 (.I0(iAdv7511Sda), .I1(oAdv7511SdaOe), .O(n8301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11460.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11461 (.I0(n8294), .I1(n8301), .O(n8302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11461.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11462 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), 
            .O(n8303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11462.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11463 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .I1(n8303), .I2(n8291), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n8304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__11463.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__11464 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .I1(n8302), .I2(n8285), .I3(n8304), .O(n8305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__11464.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__11465 (.I0(iAdv7511Sda), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n8306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11465.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11466 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I1(n8306), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n8307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf80f */ ;
    defparam LUT__11466.LUTMASK = 16'hf80f;
    EFX_LUT4 LUT__11467 (.I0(n8305), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(n8307), .O(n8308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__11467.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__11468 (.I0(n8293), .I1(n8287), .I2(n8300), .I3(n8308), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__11468.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__11469 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n8299), .O(n8309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11469.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11470 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n8310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11470.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11471 (.I0(n8309), .I1(n8310), .O(n8311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11471.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11472 (.I0(n8285), .I1(n8284), .O(n8312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11472.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11473 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(n8287), .O(n8313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11473.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11474 (.I0(n8312), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n8313), .O(n8314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11474.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11475 (.I0(n8285), .I1(n8311), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(n8314), .O(n8315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__11475.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__11476 (.I0(n8315), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I3(n8313), .O(ceg_net1335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd755 */ ;
    defparam LUT__11476.LUTMASK = 16'hd755;
    EFX_LUT4 LUT__11477 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(n8301), .O(n8316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__11477.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__11478 (.I0(n8306), .I1(n8287), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n8317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0b */ ;
    defparam LUT__11478.LUTMASK = 16'h0c0b;
    EFX_LUT4 LUT__11479 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(n8316), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I3(n8317), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__11479.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__11480 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n8284), .I2(n8285), .I3(n8313), .O(ceg_net566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__11480.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__11481 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n8295), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n8318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__11481.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__11482 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(n8312), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I3(n8287), .O(n8319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb0f */ ;
    defparam LUT__11482.LUTMASK = 16'hfb0f;
    EFX_LUT4 LUT__11483 (.I0(n8318), .I1(n8319), .O(ceg_net1400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11483.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11484 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11484.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11485 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I1(n8303), .I2(n8285), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n8320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__11485.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__11486 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n8321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11486.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11487 (.I0(n8301), .I1(n8294), .I2(n8321), .O(n8322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11487.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11488 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n8323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11488.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11489 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n8324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfd40 */ ;
    defparam LUT__11489.LUTMASK = 16'hfd40;
    EFX_LUT4 LUT__11490 (.I0(n8322), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] ), 
            .I2(n8323), .I3(n8324), .O(n8325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__11490.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__11491 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[0] ), 
            .I1(n8320), .I2(n8309), .I3(n8325), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__11491.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__11492 (.I0(n8285), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .O(n8326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__11492.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__11493 (.I0(n8303), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n8285), .I3(n8310), .O(n8327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__11493.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__11494 (.I0(n8327), .I1(n8326), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(ceg_net1463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__11494.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__11499 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), .I2(n8306), 
            .I3(n8323), .O(n8330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__11499.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__11500 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(n8301), .I2(n8294), .I3(n8285), .O(n8331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__11500.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__11501 (.I0(n8285), .I1(iAdv7511Sda), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(n8297), .O(n8332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__11501.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__11502 (.I0(n8331), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n8332), .I3(n8299), .O(n8333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__11502.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__11503 (.I0(n8302), .I1(n8285), .I2(n8323), .I3(n8321), 
            .O(n8334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__11503.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__11504 (.I0(n8287), .I1(n8285), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n8335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd700 */ ;
    defparam LUT__11504.LUTMASK = 16'hd700;
    EFX_LUT4 LUT__11505 (.I0(n8330), .I1(n8333), .I2(n8334), .I3(n8335), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11505.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11506 (.I0(n8285), .I1(n8311), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(ceg_net566), .O(ceg_net1361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__11506.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__11507 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_2P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n8299), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11507.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11508 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_m_en_1P ), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .O(n8336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__11508.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__11509 (.I0(n8332), .I1(n8285), .I2(n8336), .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__11509.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__11510 (.I0(n8287), .I1(n8323), .O(ceg_net616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11510.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11511 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(n8288), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11511.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11512 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(n8288), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__11512.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__11513 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] ), 
            .O(n8337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__11513.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__11514 (.I0(n8337), .I1(n8288), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11514.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11515 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[3] ), 
            .O(n8338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11515.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11516 (.I0(n8338), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(n8288), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11516.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11517 (.I0(n8338), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I3(n8288), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__11517.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__11518 (.I0(n8338), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] ), 
            .O(n8339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f */ ;
    defparam LUT__11518.LUTMASK = 16'h807f;
    EFX_LUT4 LUT__11519 (.I0(n8339), .I1(n8288), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11519.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11520 (.I0(n8338), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[5] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[6] ), 
            .O(n8340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11520.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11521 (.I0(n8340), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_i2c_clk_1P[7] ), 
            .I2(n8288), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11521.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11535 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .I2(n8289), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11535.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11536 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_bit_cnt_1P[2] ), 
            .I3(n8289), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__11536.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__11537 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11537.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11538 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11538.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11539 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11539.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11540 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11540.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11541 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11541.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11542 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11542.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11543 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11543.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11544 (.I0(n8285), .I1(iAdv7511Sda), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n8346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__11544.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__11545 (.I0(n8322), .I1(n8346), .O(n8347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11545.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11546 (.I0(n8322), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] ), 
            .I3(n8346), .O(n8348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__11546.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__11547 (.I0(n8347), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I2(n8348), .O(n8349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__11547.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__11548 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .O(n8350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7 */ ;
    defparam LUT__11548.LUTMASK = 16'he7e7;
    EFX_LUT4 LUT__11549 (.I0(n8350), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .O(n8351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11549.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11550 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[0] ), 
            .I2(n8320), .I3(n8309), .O(n8352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__11550.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__11551 (.I0(n8349), .I1(n8323), .I2(n8351), .I3(n8352), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__11551.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__11552 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .I2(n8320), .O(n8353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__11552.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__11553 (.I0(n8346), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[2] ), 
            .I3(n8322), .O(n8354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__11553.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__11554 (.I0(n8354), .I1(n8323), .I2(n8353), .I3(n8309), 
            .O(n8355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__11554.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__11555 (.I0(n8350), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .I2(n8355), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__11555.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__11556 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .I2(n8320), .O(n8356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__11556.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__11557 (.I0(n8346), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[3] ), 
            .I3(n8322), .O(n8357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__11557.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__11558 (.I0(n8357), .I1(n8323), .I2(n8356), .I3(n8309), 
            .O(n8358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__11558.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__11559 (.I0(n8350), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .I2(n8358), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__11559.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__11560 (.I0(n8322), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] ), 
            .I3(n8346), .O(n8359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__11560.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__11561 (.I0(n8347), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .I2(n8359), .O(n8360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__11561.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__11562 (.I0(n8350), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .O(n8361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11562.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11563 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[4] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[3] ), 
            .I2(n8320), .I3(n8309), .O(n8362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__11563.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__11564 (.I0(n8360), .I1(n8323), .I2(n8361), .I3(n8362), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__11564.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__11565 (.I0(n8322), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] ), 
            .I3(n8346), .O(n8363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__11565.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__11566 (.I0(n8347), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .I2(n8363), .O(n8364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__11566.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__11567 (.I0(n8350), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .O(n8365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11567.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11568 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[5] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[4] ), 
            .I2(n8320), .I3(n8309), .O(n8366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__11568.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__11569 (.I0(n8364), .I1(n8323), .I2(n8365), .I3(n8366), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__11569.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__11570 (.I0(n8322), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_addr_1P[0] ), 
            .I3(n8346), .O(n8367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__11570.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__11571 (.I0(n8347), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .I2(n8367), .O(n8368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__11571.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__11572 (.I0(n8350), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .O(n8369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11572.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11573 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[6] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[5] ), 
            .I2(n8320), .I3(n8309), .O(n8370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__11573.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__11574 (.I0(n8368), .I1(n8323), .I2(n8369), .I3(n8370), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__11574.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__11575 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .I2(n8320), .O(n8371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__11575.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__11576 (.I0(n8346), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wdata_1P[7] ), 
            .I3(n8322), .O(n8372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__11576.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__11577 (.I0(n8372), .I1(n8323), .I2(n8371), .I3(n8309), 
            .O(n8373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__11577.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__11578 (.I0(n8350), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_wsr_1P[7] ), 
            .I2(n8373), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__11578.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__11586 (.I0(n8285), .I1(n8301), .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n8374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5f03 */ ;
    defparam LUT__11586.LUTMASK = 16'h5f03;
    EFX_LUT4 LUT__11587 (.I0(n8290), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(n8374), .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3001 */ ;
    defparam LUT__11587.LUTMASK = 16'h3001;
    EFX_LUT4 LUT__11588 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[2] ), 
            .O(n8375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe4f */ ;
    defparam LUT__11588.LUTMASK = 16'hfe4f;
    EFX_LUT4 LUT__11589 (.I0(n8285), .I1(n8375), .O(n8376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11589.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11590 (.I0(n8310), .I1(n8376), .I2(ceg_net566), .O(ceg_net1471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__11590.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__11591 (.I0(n8323), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n8377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11591.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11592 (.I0(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/r_m_en_re_1P ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(n8303), .O(n8378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11592.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11593 (.I0(n8378), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(n8285), .I3(n8299), .O(n8379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__11593.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__11594 (.I0(n8316), .I1(n8379), .I2(n8377), .I3(n8303), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__11594.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__11595 (.I0(n8314), .I1(n8334), .I2(n8376), .O(ceg_net1480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfefe */ ;
    defparam LUT__11595.LUTMASK = 16'hfefe;
    EFX_LUT4 LUT__11596 (.I0(n8285), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I3(n8299), .O(n8380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__11596.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__11597 (.I0(n8303), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[0] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[1] ), 
            .O(n8381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11597.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11598 (.I0(n8285), .I1(\MVideoPostProcess/inst_adv7511_config/inst_i2c/o_dbg_i2c_state[3] ), 
            .I2(n8381), .O(n8382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__11598.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__11599 (.I0(n8382), .I1(ceg_net616), .I2(n8378), .I3(n8380), 
            .O(\MVideoPostProcess/inst_adv7511_config/inst_i2c/genblk1.inst_i2c_standard/n826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__11599.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__11600 (.I0(n8295), .I1(n8321), .I2(n8299), .I3(n8315), 
            .O(ceg_net1488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff */ ;
    defparam LUT__11600.LUTMASK = 16'h40ff;
    EFX_LUT4 LUT__11601 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .O(n8383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11601.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11602 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[1] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), .O(n8384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11602.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11603 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), 
            .I1(n8384), .O(n8385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11603.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11604 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[7] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[8] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[9] ), 
            .O(n8386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__11604.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__11605 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I3(n8386), .O(n8387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11605.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11606 (.I0(n8385), .I1(n8383), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .I3(n8387), .O(\MVideoPostProcess/mVideoTimingGen/qVrange )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__11606.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__11607 (.I0(\MVideoPostProcess/inst_adv7511_config/r_byte_cnt_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_reg_cnt_1P[0] ), 
            .O(n8388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11607.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11608 (.I0(n8388), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11608.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11609 (.I0(n8388), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__11609.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__11610 (.I0(n8388), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[3] ), .O(n8389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11610.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11611 (.I0(n8389), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n249 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11611.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11612 (.I0(n8389), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[4] ), 
            .O(n8390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11612.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11613 (.I0(n8390), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11613.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11614 (.I0(n8390), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__11614.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__11615 (.I0(n8390), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), .O(n8391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11615.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11616 (.I0(n8391), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11616.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11617 (.I0(n8390), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[6] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[7] ), 
            .O(n8392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11617.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11618 (.I0(n8392), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n245 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11618.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11619 (.I0(n8392), .I1(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_addr_1P[9] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__11619.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__11620 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11620.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11621 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[1] ), 
            .O(n8393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11621.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11622 (.I0(n8393), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11622.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11623 (.I0(n8393), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11623.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11624 (.I0(n8393), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11624.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11625 (.I0(n8393), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[3] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[4] ), 
            .O(n8394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11625.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11626 (.I0(n8394), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11626.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11627 (.I0(n8394), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11627.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11628 (.I0(n8394), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11628.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11629 (.I0(n8394), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[6] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[7] ), 
            .O(n8395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11629.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11630 (.I0(n8395), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11630.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11631 (.I0(n8395), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11631.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11632 (.I0(n8395), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] ), 
            .O(n8396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11632.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11633 (.I0(n8396), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11633.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11634 (.I0(n8396), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11634.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11635 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[8] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[9] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[10] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[11] ), 
            .O(n8397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11635.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11636 (.I0(n8395), .I1(n8397), .O(n8398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11636.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11637 (.I0(n8398), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11637.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11638 (.I0(n8398), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11638.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11639 (.I0(n8398), .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11639.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11640 (.I0(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[13] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[14] ), 
            .O(n8399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11640.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11641 (.I0(n8398), .I1(n8399), .I2(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[12] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_clk_div_1P[15] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11641.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11642 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .O(\MVideoPostProcess/inst_adv7511_config/n780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11642.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11643 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11643.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11644 (.I0(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[0] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[1] ), .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[2] ), 
            .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[3] ), .O(\MVideoPostProcess/inst_adv7511_config/n790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11644.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11645 (.I0(n8280), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11645.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11646 (.I0(n8280), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .O(\MVideoPostProcess/inst_adv7511_config/n800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11646.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11647 (.I0(n8280), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[5] ), .I3(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[6] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11647.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11648 (.I0(n8281), .I1(\MVideoPostProcess/inst_adv7511_config/r_ms_dly_1P[7] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11648.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11649 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[1] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[1] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11649.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11650 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[2] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[2] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11650.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11651 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[3] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[3] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11651.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11652 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[4] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[4] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11652.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11653 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[5] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[5] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11653.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11654 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[6] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[6] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11654.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11655 (.I0(\MVideoPostProcess/inst_adv7511_config/r_opn008_reg[7] ), 
            .I1(\MVideoPostProcess/inst_adv7511_config/w_opn008_reg[7] ), 
            .I2(\MVideoPostProcess/inst_adv7511_config/r_i2c_config_state_1P[0] ), 
            .O(\MVideoPostProcess/inst_adv7511_config/n270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11655.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11656 (.I0(n8387), .I1(n8385), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[2] ), 
            .O(n8400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11656.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11657 (.I0(n8400), .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[0] ), 
            .O(\MVideoPostProcess/mVideoTimingGen/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11657.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11658 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), .O(n8401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11658.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11659 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I3(n8401), .O(n8402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11659.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11660 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[0] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[1] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .O(n8093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11660.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11661 (.I0(n8402), .I1(n8093), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), .O(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__11661.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__11662 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[4] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[5] ), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[3] ), 
            .I3(n8386), .O(n8403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__11662.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__11663 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[8] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[9] ), 
            .I3(\MVideoPostProcess/mVideoTimingGen/rHpos[10] ), .O(n8404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11663.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11664 (.I0(n8404), .I1(\MVideoPostProcess/mVideoTimingGen/rVpos[11] ), 
            .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), .O(n8405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__11664.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__11665 (.I0(\MVideoPostProcess/mVideoTimingGen/rVpos[6] ), 
            .I1(n8403), .I2(\MVideoPostProcess/mVideoTimingGen/rVpos[10] ), 
            .I3(n8405), .O(\MVideoPostProcess/mVideoTimingGen/qVde )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__11665.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__11666 (.I0(\MVideoPostProcess/rVtgRST[2] ), .I1(\MVideoPostProcess/mVideoTimingGen/equal_12/n23 ), 
            .O(\MVideoPostProcess/mVideoTimingGen/n267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11666.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11667 (.I0(\MVideoPostProcess/mVideoTimingGen/dff_11/i4_pre ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 ), .O(\MVideoPostProcess/mVideoTimingGen/rHSync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11667.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11668 (.I0(n8400), .I1(n489), .O(\MVideoPostProcess/mVideoTimingGen/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11668.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11669 (.I0(n8400), .I1(n2919), .O(\MVideoPostProcess/mVideoTimingGen/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11669.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11670 (.I0(n8400), .I1(n2913), .O(\MVideoPostProcess/mVideoTimingGen/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11670.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11671 (.I0(n8400), .I1(n2911), .O(\MVideoPostProcess/mVideoTimingGen/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11671.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11672 (.I0(n8400), .I1(n2903), .O(\MVideoPostProcess/mVideoTimingGen/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11672.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11673 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[3] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[5] ), 
            .I3(n8404), .O(n8406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__11673.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__11674 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[2] ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/rHpos[4] ), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[7] ), 
            .I3(n8402), .O(n8407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11674.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11675 (.I0(\MVideoPostProcess/mVideoTimingGen/rHpos[11] ), 
            .I1(n8406), .I2(\MVideoPostProcess/mVideoTimingGen/rHpos[6] ), 
            .I3(n8407), .O(\MVideoPostProcess/mVideoTimingGen/qHrange )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;
    defparam LUT__11675.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__11676 (.I0(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_pre ), 
            .I1(\MVideoPostProcess/mVideoTimingGen/dff_27/i4_rst_3 ), .O(\MVideoPostProcess/mVideoTimingGen/rVSync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11676.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11677 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .O(n8408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11677.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11678 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n8409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11678.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11679 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[10] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n8410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11679.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11680 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n8411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11680.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11681 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(n8410), .I3(n8411), .O(n8412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__11681.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__11682 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[7] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n8413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11682.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11683 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[9] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n8414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11683.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11684 (.I0(n8414), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I3(n8413), .O(n8415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100 */ ;
    defparam LUT__11684.LUTMASK = 16'h4100;
    EFX_LUT4 LUT__11685 (.I0(n8412), .I1(n8415), .O(n8416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11685.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11686 (.I0(n8409), .I1(n8416), .I2(n8408), .I3(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__11686.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__11687 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(n8417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11687.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11688 (.I0(n8417), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n8418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11688.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11689 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I1(n8414), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I3(n8418), .O(n8419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde */ ;
    defparam LUT__11689.LUTMASK = 16'hbdde;
    EFX_LUT4 LUT__11690 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[8] ), 
            .I1(n8414), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .I3(n8410), .O(n8420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc8bf */ ;
    defparam LUT__11690.LUTMASK = 16'hc8bf;
    EFX_LUT4 LUT__11691 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[0] ), 
            .O(n8421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__11691.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__11692 (.I0(n8421), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[2] ), 
            .O(n8422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__11692.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__11693 (.I0(n8422), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[3] ), 
            .O(n8423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__11693.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__11694 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[6] ), 
            .I1(n8413), .I2(n8417), .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n8424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__11694.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__11695 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rRA[5] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n8425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d */ ;
    defparam LUT__11695.LUTMASK = 16'heb7d;
    EFX_LUT4 LUT__11696 (.I0(n8424), .I1(n8425), .I2(n8416), .I3(n8423), 
            .O(n8426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__11696.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__11697 (.I0(n8420), .I1(n8419), .I2(n8423), .I3(n8426), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/qFullAllmost )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__11697.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__11698 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11698.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11699 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11699.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11700 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11700.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11701 (.I0(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[0] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .O(n8427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11701.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11702 (.I0(n8427), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11702.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11703 (.I0(n8427), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11703.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11704 (.I0(n8417), .I1(n8427), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11704.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11705 (.I0(n8417), .I1(n8427), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11705.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11706 (.I0(n8418), .I1(n8427), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11706.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11707 (.I0(n8418), .I1(n8427), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11707.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11708 (.I0(n8418), .I1(n8427), .I2(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n8428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11708.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11709 (.I0(n8428), .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/n478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11709.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11710 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n8429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11710.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11711 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[4] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n8430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11711.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11712 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n8431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11712.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11713 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n8432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11713.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11714 (.I0(n8429), .I1(n8430), .I2(n8431), .I3(n8432), 
            .O(n8433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11714.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11715 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n8434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11715.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11716 (.I0(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(n8434), .O(n8435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__11716.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__11717 (.I0(n8435), .I1(n8433), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[1].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__11717.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__11718 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n8436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11718.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11719 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[6] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[8] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .O(n8437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11719.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11720 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n8438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11720.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11721 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n8439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11721.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11722 (.I0(n8436), .I1(n8437), .I2(n8438), .I3(n8439), 
            .O(n8440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11722.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11723 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n8441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11723.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11724 (.I0(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(n8441), .O(n8442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__11724.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__11725 (.I0(n8442), .I1(n8440), .I2(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[2].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__11725.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__11726 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[3] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[3] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[9] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[9] ), 
            .O(n8443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11726.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11727 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[8] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[8] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[10] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[10] ), 
            .O(n8444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11727.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11728 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[2] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[2] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[7] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[7] ), 
            .O(n8445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11728.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11729 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[0] ), 
            .I1(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rWA[0] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[4] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[4] ), 
            .O(n8446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11729.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11730 (.I0(n8443), .I1(n8444), .I2(n8445), .I3(n8446), 
            .O(n8447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11730.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11731 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[1] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[1] ), 
            .I2(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[6] ), 
            .I3(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[6] ), 
            .O(n8448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11731.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11732 (.I0(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/rRA[5] ), 
            .I1(\MVideoPostProcess/genblk1[0].mVideoDualClkFIFO/rWA[5] ), 
            .I2(n8447), .I3(n8448), .O(n8449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__11732.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__11733 (.I0(n8449), .I1(\MVideoPostProcess/wVgaGenFDe ), 
            .O(\MVideoPostProcess/genblk1[3].mVideoDualClkFIFO/qRE )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11733.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11734 (.I0(\genblk1.genblk1[0].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[0].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__11734.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__11735 (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0] ), 
            .I1(n655), .I2(n678), .O(n8022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11735.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11736 (.I0(n2834), .I1(n2832), .I2(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5_q ), 
            .I3(n2836), .O(n8450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11736.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11737 (.I0(n2828), .I1(n2826), .I2(n2824), .I3(n2823), 
            .O(n8451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11737.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11738 (.I0(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2_q ), 
            .I1(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1_q ), 
            .I2(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[3] ), .I3(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[7] ), 
            .O(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__11738.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__11739 (.I0(\genblk1.genblk1[1].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[1].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[1].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[1].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__11739.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__11740 (.I0(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[1].mPulseGenerator/equal_12/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11740.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11741 (.I0(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[1].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[1].mPulseGenerator/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11741.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11742 (.I0(\genblk1.genblk1[3].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[3].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[3].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[3].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__11742.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__11743 (.I0(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[3].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[3].mPulseGenerator/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11743.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11744 (.I0(\genblk1.genblk1[4].mPulseGenerator/rSft[2] ), 
            .I1(\genblk1.genblk1[4].mPulseGenerator/rSft[1] ), .I2(\genblk1.genblk1[4].mPulseGenerator/rSft[0] ), 
            .O(\genblk1.genblk1[4].mPulseGenerator/equal_6/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf */ ;
    defparam LUT__11744.LUTMASK = 16'hbfbf;
    EFX_LUT4 LUT__11745 (.I0(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[0] ), 
            .I1(\genblk1.genblk1[4].mPulseGenerator/rTmpCount[1] ), .O(\genblk1.genblk1[4].mPulseGenerator/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11745.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11746 (.I0(\la0_probe3[0] ), .I1(\la0_probe3[1] ), .O(la0_probe1)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11746.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11264 (.I0(pll_inst1_LOCKED), .I1(pll_inst2_LOCKED), .O(oLed[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11264.LUTMASK = 16'h8888;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4  (.D(n678), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4 .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4 .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4 .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4 .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4 .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4 .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_4 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3  (.D(n655), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3 .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3 .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3 .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3 .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3 .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3 .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[1]~FF_frt_3 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2  (.D(n8450), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2 .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2 .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2 .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2 .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2 .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2 .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[5]~FF_frt_2 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1  (.D(n8451), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1 .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1 .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1 .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1 .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1 .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1 .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[8]~FF_frt_1 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0  (.D(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_5_q ), 
           .CE(\genblk1.genblk1[0].mPulseGenerator/equal_6/n5 ), .CLK(iFCLK), 
           .SR(\genblk1.genblk1[0].mPulseGenerator/equal_12/n23 ), .Q(\genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // D:\workspace\Efinix\Titanium\Ti180MIPI25GRxHDMIV101\src\common\MPulseGenerator.v(54)
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0 .CLK_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0 .CE_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0 .SR_POLARITY = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0 .D_POLARITY = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0 .SR_SYNC = 1'b1;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0 .SR_VALUE = 1'b0;
    defparam \genblk1.genblk1[0].mPulseGenerator/rTmpCount[0]~FF_frt_0 .SR_SYNC_PRIORITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_a648f924_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_a648f924_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_a648f924_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_a648f924_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__10_10_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__10_10_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__16_16_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__8_8_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_SRL8_a648f924_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__4_4_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__4_4_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__4_4_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__4_4_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__1_1_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM10_a648f924__2_2_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_a648f924_214
// module not written out since it is a black box. 
//

